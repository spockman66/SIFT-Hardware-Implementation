


module hme_gpio_v3 (
	  gpio_pulldown,
	  gpio_pullup,
	  gpio_intr,
	  gpio_oe,
	  gpio_out,
	  paddr,
	  penable,
	  prdata,
	  psel,
	  pwdata,
	  pwrite,
	  pclk,
	  presetn,
	  extclk,
	  gpio_in
);

`pragma protect begin_protected
`pragma protect version=4
`pragma protect vendor="Hercules Microelectronics"
`pragma protect email="supports@hercules-micro.com"
`pragma protect data_method="AES128-CBC"
`pragma protect data_encode="Base64"
`pragma protect key_method="RSA"
`pragma protect key_encode="Base64"
`pragma protect data_line_size=96
`pragma protect key_block
T6mSsLy2Uv05EC2MGLuDqqu25GzVpLwjXHOwMnwmXysbGfOqgsPY4yjmFCxo3Xs7bJD1D0Sw21fl1w9wdlvTfH5pTXmgxRmgrhH+oWpicMfOrV68w1uqUXNpoNgtykR6k6OqfX10EBJm4r8z1eUj80JEfItOZHjvdUmcl+fPvE8=
`pragma protect data_block
ackkGUSoYe0pS9luGs/vkiEY55w8eLD3Uywt0l/xL+uZV/CRPZSDYjX4kmL+bLX6o/YuXadnouX0WMNfF1OgWqwZ8m9HSO4DDISxBlvzpu5+mGZK9qqCi/xokH6xDdf9
+qeluZ55hA2UXPiafcQEVQUu89IEzcngSXDnSaM7JSMQTndY3L8/JN4LzBoBsGPySeVIJUZzZdzZCjEXsM4+dvyntqkVExocQeE4WUphAnT8noIqiwsAFZmrUCOGDpUe
sh2u0s0vnSYTSSyRAfWAvbe/rUSg5EG6nicAOvLI1hXKiCbRJr2HgYyrX3ljAm2IgXg2XmkZ4vgmw4SM6tPTg5v9HbfcPmFUUmo08cXfxIXcwkmqBNzgOWFyC+bHHC9t
HQ87wozU++4tjaY5ADzpvIsRwR1grmKRfjQOnCK9SCrM+kN27h8FAFeHuGV32yHwjPHRnSI97ITL0HPkBzCDWB0PO8KM1PvuLY2mOQA86bxWF0NkcwaCqp5lxFQaBPz2
a45AQE+CvRbtELf1zPnpol2v8b+1CDktX25OvW0ZSMIdDzvCjNT77i2NpjkAPOm8oCnkYLAiWTkxH6VgoGfqfTs+FcowHIPWZY/nMBcBQ16jUIvDHlQV/Yf1TZTya4W/
2RXf2pgu2MXqbGQ6OE0BbFEeXccT4DGreDvm6Z4qKkLJmWOLmwP80TzofK7kt5ggzYl40fZuPBBOdfuVHGnrg7NFPo++mxCzlvQqpmwbIvlKpACPfvP07+XEmZDSheuq
dV8AIa6MqgEIed6XGMKlJUZElKNnIQjB1P1PJnXGVnN5D591m1DEhvDVybG3WfaV9sJb8XraXyd1HU/q+2+hT7K2s51uCbE9Ijxyu6/hdhlxDUrWHaZkCwZYKD5WgVE9
zqJMqBnyV8VNXWHPjDM9ngdew2bQpHOMFqaqCa3odlbu67P8cI10Z7DVSmpQCOCau7KjAfW8bkIYleZe2KVNvsqIJtEmvYeBjKtfeWMCbYgNR714E4BStABFikAVhWf8
cEi3NiTXa6JVv7kzhOq/iu3+jOI24fOkNNF7yxZHt4JfL4i8gidCQA7qCW/D9P2aGKhpguf+W/+LZY8pZkI0Nz0KRX+KNmxhfew9TwEGn7dO3SgAx9xfoiAnyY0+4Pxs
XGmVy2AccdP4MESvhZt9MXeeRNUN0/8ErftvPMxlCwqmcpwpF3ppBP8M4gl07I32iu9v22qVGap4R7Tvk0R3k2I7dvVMBcjUzyTyZLroCMy1uz/HWfaVk45A4w5WCgOh
ScVQvk8DMO5DDuF9FF2pUguWuNWGFOJJmzj8GKXb+jT7QubC3/TT27nbnBh2r660ryUSIyogEytZ6e0n0C6t5jgqKcK8Sla4KV2Y2I1W+ydMmVNP1BIGf6xY53a85TVM
/Gs5P/LZJbE9KhZcZlkfET94MVrMJMYS8gkuM7D8CJE6QXvfzuwAkWkcEmuKcpwXgWkQduZb0YEJnYaOMod92j8hKOhYfOrsTed6FyIj9J1zT3gw84We863umFpuW5pk
+PVBEc4HGKqnWtY6r+M/PNvCWB80E19SN38qds04zSYDWCwdKZeiBhLVssUtd65sNP0JiQkXo1yDxmlna1c84q9CSW857753uy3+8TtuanIoqFD0mSSjK4L9Dh1EsHFM
zny3smSN2QztFV9NT/Df2kNTqhHgSCWEBHbvphiXJUOGbZ3qb9/l4p6WW3t7fLbZ7LcCRmk6nR6jIOGLVdltjCa0FEfXheAFAizHVYq70hspIOlqF4YjsUGYX9FksDlJ
4n/qKMG9oTrYHs2CHemo22w42lE1AMOVfz8g4vWxwK1CkT7tAAOgUXJlT5VwPfoE3K1fOBZZnlfOfIBJc0yqGHlfbErMRjQbIh2q9jBFWwomsM6jX4L48kWAOwAUXu9D
jMk66Q9hGTyk1QhgmTXAlHna9ulUBdHArB63ndSvhZn2wlvxetpfJ3UdT+r7b6FPNT4CHjTvSnmcRkol3D0w9zjrlmeGiTQtgBIadeGWOKxAli8MDp9D9xK65ob130Rk
tqxbwyL+jBIpZPgwdzkNu/UoazOtaeoOlYdcGkpmc1OcccFLxhFi54QfWiHZ20r5aaLWw1hgA2cioJpNhrm3Ao/DNc6/1892EAhOVF0Qkutrz9tX0axyrLDGIA/ksMv6
2Sb40ZWZ6h0gqeASI0skFZgmYww8ZjJMMxt7FIJRwsgCxCrdl1t7Y/4czxGpMpB/Nrv6c8H5b8R67iAMJCpTXzEZ3KxzJQJJZw3mriBw2sMO8lSIQ9qhhuMuFsoK4gE5
jtgsHB+iz7McQXNy5tDUUGPE379Os4LyRWwJXt+tXV1kSBki/h3jf7BJE2wC4bmNxuadYM8F4rYeASwI/uuluI+AzLpLcINoSmxMDSffZifg//Owv1VIhtc8qeHbLOt9
iO9H5pN31QjslB3HdgFKNoOp6DSgU4jRcKgKNnlCsqCkj/jBhzyQkNN1dPOefjvmbABL/e+TNW2RAsiBjyMHvQtZlVP2UNTSKiMHK40RFJTba4j6vk4HPEkKQwpiHZev
rlsfX5UuQdrVLRmfWkYJpT8x5eMUZH1l0gFfBElYNwocgtdtQ+L3EMmdMEHCw08a4lgstIIz5QqpWmZSRJ01oL/rO00k/3Mg1pvDoOU3FR5GZY2LMH8D6GKeT14BTUGK
qwF+GPLERzJtauGo+jub3pEGiP7sjMbK0RDFTJGakdFrIX4rroHJLn/POlGgFJfdiaem1ukGilIt9dZOyLV69OlV6WYYqyepL4MzCmU2tNCJPwpznkmbKZqSk1sjxaSG
CeV+2OMf07h2J5aq4THtAp3ZyL2Xy/7sCdhhqdFekBwHubWLOmJD2gOEKX0XIp09Zx0t3JCUESc2sBCfgCKrTHdvEkrs5bFmCTC4jygHDIKqD6zFTwnW/cgmJHALni3N
NSJhx4vAYYfwFgkc/Vo8wEinUDbvdrgK+HlhTdAluY0T8hCQC1Sgo8YycmLPJ/XP3BVioVZKgIbUHIuO1Nhz3Cv5Wek6VtMHdDD3ceYFTaHjMH5sFmbqleJH8J4qnozj
+JqOo4hg4NKfV/r+06n9wCQj9y1Xi4GSh6P8rIIwFfCO835ey+ooYLhiqlXAwzABGP9g9BAFkteMwJL/YLIMUL3945+YdzMogyswawEsbeWnbeHNd8SGOd2CeGKf02La
Ik1wPMAKeCeed7/Keo1QyfGyBGn15YSZ0jP2o8OqS/RUb7NvbeSQO1xQlsrqXwl+Qyft7mB2jkYs233aEylccFSjJal0qe8VM2VJDv3W0u5z//pT2VvkJDUyRsohGsgs
yogm0Sa9h4GMq195YwJtiOpTvrSHMWLC7nhhHhx3BFjKiCbRJr2HgYyrX3ljAm2IGDJEl2xpu+tdbRBdK/YUaY4wUO+TxBggGcuMQEDz7mfEu2a4Y/c9B6j4FZ79wtGF
dLSnI4VoaFmT7+F8G2EMXzkgsS+9DQJIN61NZtAFqKltxU9CMoxr8dck/Uk24pdmyogm0Sa9h4GMq195YwJtiF2r3YE/WXhdNle8RMuLfLKAaei9aZAUQ0FFlWnuw08Z
yogm0Sa9h4GMq195YwJtiAJAqSWQQkeSLK++MQ4A1XhajXWitdQ0ATLvLB3QYjMAyogm0Sa9h4GMq195YwJtiCsEyR8c9gNGL2miCZpbLdWRMLUZ+N5nEeMtyBCfAqmJ
yogm0Sa9h4GMq195YwJtiAsWcQqRL1EsiiWOFG9TOKkGeGPofHoqoLlWHQTZLXtxSENTCwsafwJlrF+9Puuja8qIJtEmvYeBjKtfeWMCbYhdq92BP1l4XTZXvETLi3yy
CTaPy2pbnjZtby3pckT9OjkgsS+9DQJIN61NZtAFqKkE2kvSZIjJsls2/GQ8P86ojjBQ75PEGCAZy4xAQPPuZ9uK/gC4R6VK4sAWG4CEsO4UBO4wKEbCbYephN6fHqdS
fDiseQJoIo+bdxzoDe3uHMqIJtEmvYeBjKtfeWMCbYgUIKMXi3VnK+xXQK+bBIcN240Ztijfg1n+ndZoAduGI7SBg6tblrqP4XEHXBLu/UywTsTLuYKtDjjAdU1Xi9U7
yogm0Sa9h4GMq195YwJtiGkcfJSa6RZkImABnjO6I/0Rg1X0pA8QvxBPxLdX8XfUUTNOs2R89rziM2PXDAvDptkUkRhUpu1xxYYmXZZgJO1BCqifYFhu1WucEoYdu/p5
CcrbxEQRrfsmnDsAVGjpFzu9As58ucoYRRq60QDPcpi2qCVipODOAW4tj7A5eJOu59KZ6FSxaao+HObQ4DqjsMHFcOKmyOKC51VV9p0uVmy6Bl+3VTvaVFSgONkk/rV/
reWSsWQXXMocb3XsHTPyf4jgo1r4At7UVBuEPHXQxAvfFMzRVt/9BoOKiUMDWWqLZouw3RWMu+YvF8WAFa4S9fGGvVto6pVUQ413PFHfUN/BxXDipsjigudVVfadLlZs
gtf54Ij0qkI6lVxBPSnm7vIr/37fPkJjmAls7Avk87Eqr8lsIYwzcraSD/9hOp4hXDbxztMaYFHcdMDYpv8KvgD7BUUICKXau9cmNxVeXzqOKqvqUD8OwZZnPCToebF5
bP4j904rX6tk/s+jIGgj7FQQ20798iDc2BZ+FZBN2mpJCkmySIyWeqZW7lJig2uYDUvzOjSd64advM037mYtiknjj/+eH21xIEbvNE5jaT+OTP3Qxpke9p8I6n4qMJng
t9ubA1K4NW8HYi4GWanDaK4+lt3tuWqrJsikKNLpCaE+9WGSm69Bzp22fxa4kXJiNGiSNJH29rUEkYG9ehWjiYP0KPE83/30B8to/pTU1LSx5EhRWZkG1VewEQsLLtK7
taLoA9Z5hgvflfMp98ZG50Xo2xcli+Z+moKpbifoB5qx5EhRWZkG1VewEQsLLtK7z8IEfjs9ebG9xWm8tPxsm/WvUI18eCmCM9VkwmG6AK8WRFyV4r0ndpDUD0D1LOh7
CdctSO240Q4ku7j1ojWAUdIf96ypRt5JXXOxj5LMEBNOhvSD8CbDlqykW5SUhhqRvLXE7RKPVwI2Qok1khD+6zx3JTFadOgTPQOf1s6nAbDKiCbRJr2HgYyrX3ljAm2I
v/a/t6irYfmfU3nJ5gupifMqkMAVRS92vc9pXLDLA2QGucNBf/XbUoC1ZEberrO2lnPivBUZe/WsZLTNFQ/kfBrPfollDFfIhs6UTxAkTtJPFxK+AHpRknTbVpZTN6gg
C7yRzF1AWsbLK/RNuRxKL/odV5nCS7D+vHE32eBG8UE21edd5XN/3hBGKeSz/jQR0AJr4J5+CKrU2oTZcgcczqvETd69xBbGQ4a9M9cEdCmm4zn+OHEiNQ9Vde1c4TfL
MXSg6+ihBLPRw8Y7YYk+NMiN3B/CbnFRhO4ahUd14v8Fsv4YwAgGnrpPW45UEyWO+2XNnnxTr+jYGREIDUEY/Z6WgEDY69HcfXKpK+rkgsG5MStywM7NUuCZTTmJ0ru9
12/CbR87fuauBvgn0tRoNZAApxkSI2kp5oiY1CB3ICAp59t+wwWdId1/9jrXroHdMH7AQR9SYrlYTviYwCaYR3/mVxN3wA7nmGgUnBvYvBrJOoCE8D0nTuqbpT2enK4s
0czsatyKfMehVva3Iq9Ftlx5BVf3NDTxKB6Ga01rbvZDKoMvt4iGFaCRe4bauGnm0oGEmcvF2g26WeYqKYw8FwYIeQ3K6MvE6iMIgklc995zaUfuOEVvEGsio+OCBGAs
XdArF/Pt/dsWEv8N45p5mW2434lWojCOXqHZg7vCvBVP1aroBjHOzMsMBPwoC5rpuhcdrH3UVekyNGUQsuvdAmM/mKcDFOc1o82cIkgYeyl+7Mgy1PmSbUi2hCPFpQao
G6FDkHyQPjdHf+NT5GGId124TedTsLdB5WchrLPNwSbWY8vU0lRnc9IJ+fNW31co1YtTUdRtHkFMpysFvQXoM91hEcFnCHwQKWftsKHsn0BQ3rEHKgMMSgF5xJJMmd1u
DSwaN3NJQ7x3K5Mhla1BAwWUZL14VofUCiU7oayVNxOTdn/LDl7uJMRxBJJWQ9Ziga/Y7GcyHwkLeKtQ+hBrisRWQRmmtTt8sse7yKGLCfSDwfEJd5X+BiXNPgERjEiJ
nsT9uD2+3vQCS0uMH/h5G5QkW/96Dy5BiA47gOmxLkWF7oY+FlavaJZ1zxyDhJmgZouw3RWMu+YvF8WAFa4S9VvjyhWqYogAX0X/+7EtE2N7iPlgoJl4Yt/oLWjlQi17
OQQzCoaW5JIcKyPb7NXx9/b4U8YA0GmSPV1lDuPjQUhfcOI4278X1rkjfFYoFtWxsBvi9Us0YnCymNYXydyq9KhCwrtYGr1FhAxXLrtrtII4GJKAfo/t1P98KFpqBUGm
IWkuJ/CpavNEySOIXYikISAI4FN+piE1mAXnfLRiexf/9h5AQyNdfcO4WQPv0ifsPqFBuOLjcY3FCLGBmgVI4hlejFF3jTYuIegnwLLJ7ZGux+UECgLnHpeajnX7z3YD
MeL74aNsOEaxmxJ8YMwha7sKFbaPgfiNoS/OSNVdsY1gcyXEc47h5U1lCJvT5X5fnnv/apRMNSTZi24Q+UtSlgcUYCAthcIkaZTLC6iIsP+Qu8kvdDYEQIBqeUoLEhEW
A8Hrm6ML4ARO7OkzcvC3AY4/Md3e5qdyABFf+TKvU1NIgVlSNS+u4DwD0VzRmecZre0GHP+MPl83cJ0meDvY4pqV1L1tNMrd/sdf3rOrhV034fdHMZqt86i6ZnhxuRtr
f49k4D+JIZ/1KvG6rVQHsvQGdao658+wmtbvUxO0X/2z3/D3/hoSUFrKKdNEYpNv/dbpq0QyeVmyW1gFM+IWdU7R4ZiTvENkRZf2nEBalTqGcpTncTeK+1OwL6rRoRWx
C7nXbNZ18afvGyhCzgaYZVV40H+Gx+yS7hNaTV49p3u+d5CHFfoejeFG6SBhFj8/jXijO2IYkyxfoY0v0bkK09U8RqEUI1lB1PO+WFxkPdvgEumW9tKhqMRBssmooV2R
KQhA7sVEvkDKU0JKqlYphFsCoH/MSl1qeGOfwQW2q9BuF4B3RM3CqQaOZxae9liBc2dS9CrgFgZUsuVC9dG4h6lBQJ00pvA/S5xXPlzNW0tybna7jUcVwI6jZXFC3U8x
tUmsIdO7VrlmXE6n6+iQ1l6vhFcsu+HvuU12+P4gZ9y449zCM4RSCpK7RbY9SRu4FkIoR/RjjbW6P436KG+8F6jnE27CXHKwPP9Olb0hGm5i8T5nOtVMhYzxMThjjdbh
Gho7Z5R8D+JcT+nBsJkaaExhJy5LIv5W7lLnb6GVsJqUdbsNE7LbGw7w9Q6Xpnh9xOoNMeQoUBnZVyGPlSeaVejubtet3XddvuNvTxQhOz3GTX1SczTgi7h3Rx09Z8rI
yicpjpHSfFj40tSJDsrDJwEeAcaYnAUnEr2mqDdSFAIz145geMTO9YMxs+gz4deIDT09tdQhYGr6kH687WWI1fqwgw2SRqo//5JbUILC8CuQ1OVzIQKEN4QSS768i36y
OGyxN9TrJu+dUK15tl9uOrt4/C2sWtlbctVMD1Ku42WbUdsszNKyIG3tUtVGLnAGUYwlsalS1yHdWjrbKNmGjwbqCh2dpGHYy7nqqsTOljqGcpTncTeK+1OwL6rRoRWx
C7nXbNZ18afvGyhCzgaYZVV40H+Gx+yS7hNaTV49p3u+d5CHFfoejeFG6SBhFj8/jXijO2IYkyxfoY0v0bkK0xHwl+YShhx3n7LuP86qnnOiaJU/g41A/YpWY7VNmRhh
Rcdv4KTpZwegfXAwl6l3wyQ0dCMGfo/w/c6kqNLKgLnKcAFy5/BwO+MriOkUGoq4qIMQx/pBrhZm1bcnSeRUkX41jjarY7IvoeQvQzrXhu//e9DDKnwyK3q8A1s7U4Wm
kqpQJorI9EDwyttmu6Q4Xt/gS4Qg4pE/kZFJjBSN02/Mtp9rWq+rs+1lF0GjHaVLxgf+EU4Q9NgxONT7+rxZjHSTptCzY5aQeEZBXHVOsKFDNE3jA64bxqGdMGuQTpqO
T49rHoO5xIbPGTvXQMds4i+fX79t3xX2lYFG6QDr4Um4SsHfkULKjSSEW3JB1w74SwR/+1+9ZvTIj/iOND0e10SYPxD3wbU+fZnTrrDm+lSYKdZjTB4MlI3JnM9aqMLT
a2KoULLq6hypwk0Raj1hjVFYGc4We5T/NMjSa5FlsEKR28GJRanXsc9I+Ir/8Gqx2JkS5owtcQJCoM6OjSrddnx7b/N9zIEuHUNRc3aKeIuIer2Dk0Bx1y2RgpvTnwif
0EaB/n/unS4C6b9GFtfvMOnIk4WShFniLK+1J0/NykbTyAJGyYF6hHDRmpe3zJVFtojRPkTkXRq8h2pasPWqh6Le0W5SgqSTdJJI6NPZWcJnB6LEM9nSpPhnaBTjiHmL
Ewh3QAsR7qoln98STsOJedZbwyCerLFvdRtKobneq7ZYojP1D2/DHhHjjZNzdsmv/Y7qS4RL/TK78KzNw3YYOEiIPCvLiITGTbuemrKIfd+fBZokwhfdJQpfSPmgL+GB
ot7RblKCpJN0kkjo09lZwv1pCufZ1LFp63nikHgtp30ZdSmYNLmIPtQ8hEfYKnebRiueQ234llyeItH+BctpZ+DrjyPA/xuNBTri0pk+M6rQRgbyEoY1m2+sTPXieLqW
pbkhKTIbH8R/kv3tSH73Df970MMqfDIrerwDWztThabehBzJAJnyJk3UFIZpmcUm8taGQBJYLmo96EIMaPvZl5kr5sRrhag2TYfYYrnEM+pwz0K6j86TX/sLbB9es66j
NJFHZcJ0eFg/oQIyuqM/pLJToRMFyAtuv+YVASY49jwvB5m1/fjTPeB5j71UCY127xwF8HkY+plpsL0Pk2Dadxl1KZg0uYg+1DyER9gqd5tGK55DbfiWXJ4i0f4Fy2ln
4OuPI8D/G40FOuLSmT4zqvUA9TEyK9A6l7bHhRqkNJckXK/i7h+bRnXA7B4i/cyqSLLroSprhOQegqwvMyvP/f2Gu3CBe8VPcEM29pRInq4bVOiIkUhSfM+kKfNjW/J+
/Wio6ADOF3JwahOaOHgoX0cT2PxdgjcvRBdlodixE7iehZHCTdqrD+xCvdA1N8O8GP8Qu8o90p0AMpluc7oC2twsuMLtAyRMdS+i/36tQheMU4C9c2qtz6jfPv08IWAe
WvevqcPjqfSCR8VKAQQNF/bOunmCCjQNvda6Vub9oIPKiCbRJr2HgYyrX3ljAm2IcGa+n+5IFAe8rNxPxC8CfMqIJtEmvYeBjKtfeWMCbYjLu3YgH2HWp6OayWnRfRFD
8FQYpIn4nYH5ceHDpqhSWwVYxmETSdogZBoA+g1M7jcWP6Bthr7g5JA7Be1huf4gOSCxL70NAkg3rU1m0AWoqYkdbFb+qB7mWTHUoCffro3KiCbRJr2HgYyrX3ljAm2I
3xTSfjfxBwGljG3TplB5m8qIJtEmvYeBjKtfeWMCbYjphjn/1BABLTet5JOWZLKpyogm0Sa9h4GMq195YwJtiI5UhBoYESnv754phy64HZeOMFDvk8QYIBnLjEBA8+5n
yeNXpdQhxjuu+VVoalBKTArkSE8X/j5Jq4I2Hjxr48k5ILEvvQ0CSDetTWbQBaipAFpG8CWKExA8/61i9sMYXcqIJtEmvYeBjKtfeWMCbYivyFnwfwbTttyLomzYg3yC
89zFHaTziN1BZEhM+NF9lMqIJtEmvYeBjKtfeWMCbYgcsbTAq3Yw6LwDPBjVnnREUW4oTrfIMxIxwwwuLe7fcDkgsS+9DQJIN61NZtAFqKlcXfd6ADEj4apqMp7/HeZ5
yogm0Sa9h4GMq195YwJtiK/KidG/K+uDXdgGxDPxcb7G7+dJXIE9wP6YA21fyPWsyogm0Sa9h4GMq195YwJtiF1HAOtJgYTWXqtoqMoKlQgBZ7lTelB22h4r4iFCn+QD
yogm0Sa9h4GMq195YwJtiK2dM4Daxdra71kSImyPy8HemEdvKpqX4icUe37ydUX+yogm0Sa9h4GMq195YwJtiLpmEcc4fhWmjsQ8N9sycpLKiCbRJr2HgYyrX3ljAm2I
dIR3HwIGiasb6/4RUKeIbcqIJtEmvYeBjKtfeWMCbYiUH4XRZsX4NZpTUkkMt6Afyogm0Sa9h4GMq195YwJtiPdasi4qdDCciEbiBSAz8LqXLbZOVik2e7HxsdW0ICzr
yogm0Sa9h4GMq195YwJtiCavaWAfvsxYNVhmy+7gUybKiCbRJr2HgYyrX3ljAm2IgLmVOEg/WTuvJJQXSZITPZ0yUkZObAJnqumXZHwGLIawTsTLuYKtDjjAdU1Xi9U7
yogm0Sa9h4GMq195YwJtiOCl5jCNrFA+7N6UjejQaOrKiCbRJr2HgYyrX3ljAm2Ixb7HlRlHAw0pxWxs0kytGI4wUO+TxBggGcuMQEDz7mdHayaJSDEGOEFMHhYjFbjs
WSQIiqA+WYjdUvl/9UCkykVj4HV5OsPQqRZYU097eP5wxnwMXi5n2fsPPWWepfCud6DIp7R+hJYyz6SWoNIFUaGBkcT8SW3ROu2VKcHuv8bbECuRCYtbDrtQr7MyJepw
zcSu86t4tnyUJzt55pORR5EaQ5tXkTpkgUfUhp5UP+90xwe1lyMP9kBqgYv7/zGfDCzpsQ/p0z/uF3/e7mvbK0GhfI0M1D5dMU31F1CY16sUwpGyR7R1M61+P0geG2MH
o9aBMDecSw0yH3jI6hz3g04gMvV3VHtk8w1o2VX5IUMaAl0UKKH7VHJzaXYsc4RUO7okkiocwh8WXf/ZRdMnsHNdRZ6BUSL+TNEml1LbmVTutHaH0gYOUFf3OQhaYW3+
RcuLYCkJXgHZU/pkXy3Jqfq2XAl4WtgphA9gBC1BthdFAeOenVCc7n2F65528VV23Rw+LGVJxg2YUdyECPRs5TOpktyPr6UKSFVxhUjI9OJUMWVvzW3/UnkLVIdR3+eh
RcMX0MUuwDRlyAVIVB0ioQz95d3a2zj5LqvzLM38viI70iyxxFo7/3WDmqphdgGUYntmL4wjwvZT8eTsgt/OKjehNV4IjZc/Z0ZgFXXlftjM3v5jDkxLybP0F2N1ywfc
PFz7I+MtrMxel0KTvZ6hDbIYngxmBvSoTuK583z3rvcxmWqlu1aYk7QlpqTYBOLrry0kuMkxv2hWuS1/zVJTbVNl3exgn3Et3AdFXsIWfVtbGZh9O3t0qM7jUCE7dzUt
RcMX0MUuwDRlyAVIVB0ioejZSPvp0s3rxmh4H6PUarC2Swj5ZmcMQm4apgWixqBqGzSsTeMdAcHnoL6QH9KDTH6YZkr2qoKL/GiQfrEN1/2tQAmeUqrZvVXk0hx+xHHv
3Rw+LGVJxg2YUdyECPRs5Vo1hEmvg9Td2ePhWVzjamBcXrEOI2gz8mSDj4T60iBgeUbu9ASFj23PltIMgUR8YsiMwRadfkQ0hEjdsYh6PzjHaubgsYGjyz9m9KAYHftt
EIFvi5DCEmww3d+4GZ3YuQ4qesU0gOozK+00INldTp6G4LA9CRkT5tcnd4M5acAdKc7FE3NzJwbpF6rWIo2/4Yjt6F41C/VBpfdA5iY7hSrPiXeSu0eDhpfE7KIItCL5
pGpzjX4hv8luDiW8ph4+WJ3Sizr6JqgOxlfxeGSbNWCLiZWhmigcjIFDWkLdsfDduJ7/9jbT0Wjl/dT+EO2cysJ4aVU78MKCa/37RhMQ4hPOGXKCMhJ4sdyLcY+I5OFv
OSCxL70NAkg3rU1m0AWoqX3myUWZkgIUdk8dBQhVPKPKiCbRJr2HgYyrX3ljAm2Inx/QzSexDR8XPcE8ZQ5jgkdsTxHSMe8UaREA9s/I8YFAXa/+2bFYEaVD9WuVNeru
kN1PatxQLn6ARD8GGEf79T/ZLMjBq/Lv/GR4DQlCjnLqVauzqxLm1iJvhnD6aFxTtNH00CejeTRyTaSa2BH+/n9LWgEB/E/Xkp31z99QYRadMlJGTmwCZ6rpl2R8BiyG
VsJcvdegHYpLEvsbohj/tt7YN+iWSI0zfA+1UPUf1bKGVjqmFZ39Ht51HqSqfRVpRtkv5oPUN0pWdD3TY2HL9Tweq19nu1vG9NZUbgtd09LyGfdepISTmeLzOiM2kUV8
pI0Kk+EEZYSvX1B33O+BFE5qh3XK7ggPckSWQR2advGtlj5d1KQfiVjqiZJJY1NX1xddRxoNs2sCZsMiA+rwIGFAy6yzdSNlD4O3cd7q1udHbE8R0jHvFGkRAPbPyPGB
FDOMdRbHGMMeppnGMSne9mFAy6yzdSNlD4O3cd7q1ucgrrXNOh8NtY/+96OoEPelzEKNmfsOqmS3MBDw3qRUVv1Zw95pNj3JZFu95+eISkGtlj5d1KQfiVjqiZJJY1NX
achWMHOY4ATRGR2cTXFmM6ZaWqNwc0chdRqugeOHo4mQ3U9q3FAufoBEPwYYR/v1hhIGTIBWmqL2dH0nH05MhBrUuxKVQwhUCtprYOFkth+00fTQJ6N5NHJNpJrYEf7+
VZFleF4JOPCe2VGU548nNzkgsS+9DQJIN61NZtAFqKm5F61Rp6mcnK0H8vxKXEuP6eNT9y27+zjQjZmWb50EZgz04S4OxN/OcZBeYHibMdsbM5SiojCpJGloAFhDbJSU
INCuVEyqZcG2ohdbPNO4pRszlKKiMKkkaWgAWENslJQ03jhyVi4aax77/hDaecKQvA/0ID4wmCHqahac95c/YEL7pb/ODO7F/qNz/E/Bf0UeVXDS08/1+MFN9qcHIjeq
MWqm2gHqZNrhPiP+ElthfE0KNXlgFaRzw1gfyBbvLnqTIQfFoonjtjEJUaYwE5DWmcze43Cy96g/CGZRE3IcVx0bIugvBpgojCdfS5uz9LCFUz44kvW1xmlX2a/Nij91
XMgdnoLxMDIeWhjqBZfS/DGZaqW7VpiTtCWmpNgE4uvd4/TZcqyvI2uPy8GyiyJjs6RXVvyDWlnrDg5qdWXL2oI2lFmzDgoIHcMcNr/F9Jn6HT4JSfSGlP09vUJhFaCz
PKWlR0hjhtx1yuJ6Q21q6NcXHf0MHniXJt0CGDmUT7zutHaH0gYOUFf3OQhaYW3+ClguhGcJ+4bGoLjU6vV1xtfp8UpWglmBxgiicfF5VY+3dHAXdg5TbnlTuBdf29y+
hzWVhFDajcVe8XKvPpRmpYGB+mfoLl4wAyuVC+qLUqTKjw3QWI7dFB2Y3BjEoINWkyEHxaKJ47YxCVGmMBOQ1hSINb/zIZIPSazMHT/SYnptjZZwnJ744AArgK8RB4zE
JRfl2WjrlSNczxt5OxxfOoGfBrdsnqjaYO9fRagm1WZfwiVu9GXTVRHYOwgOgQcdf3iKdJAaqEPKEbJras6ZryKBVdptBe0/8OubhaQSIdP13WsoQBVOoaYKRA5BH2QG
/n/dR59HzsrH/CcLXVBIqIqFWa2DAEn7lQtw3ils7mFr6Wuk4lWARKt1pkHynPowEX6N5Mz2NWrbiwz5zVoijfsUkrZlgVjhKXMV+myXZJ23VZuTB0sRl3rV4sPuxwCx
MpJZUv4Bvu5Kjj++5WodqXPzj//P1Ujz1GDFMQ+R26MoM7cKiha77j2c3B9vxz4/T8O2Idv5Lty6Iw3N1D32yvKYNEm3ijM/5s7S/C99s2DEeI75gEf78E3VrWh2JkwD
lrEyoyXkxTErqHpThIMXBYeW4pCn3/lYCeLqP2pC4cs2iDCYta0llQdYbiQVTwjWFwUs2Ji+U++FT5930pMWPYQVh7xbVbuBFefH55p2ni4r9MNaHgr1voc5tGXpPjjH
YE76ntUVA50ovvYICcsq8eBKCpdsx0HR9sRtlz5mtMT/x711Ge9Epw62zsecGwLFQaWFbUG2VXwri8sg1g0pQ+OrpJLi4CJl6I/xKvtnEVWo3CNEkwrMz9Al8FtpnZgL
CTwx5qArtxawaiAJ43HyaAgoTqo8t1b8nIIsWVe/SAKcD8iPmzDAjWrfnyvvhyC9/B73t4XnF2ITklrMzn1RUfTXQrr0rG7BC9hdj8cNrWgPDjNfmHMmTxkQ7Ryx+cFN
uKWycJwZqY0b7m0VJhswFqTNMAt7mqEgFUalHJyq1cjdiiojpG+oMb1HHhf71+BaGuQp0mfb9PAzRuYtgc+U6q8TRTXm3+yE7TFu2IFluzRDGY4H7NpiBgRd8sjDRSqG
8CUmRND0Gp0tStOB2EZlmBtvr49b5sCdBmSrKlvzfv8TaSqWAYoSKtBgI/gW/d7XZJLq93ZvCDX8VAWmTSAJj+FlkhIYlQwpXHTBw9VxDVNoauAIg9Qa1wfjgGmW2NqT
r2+gl7fsrOi5Txa6kpuMJnZToiLMIqE/+sZWZwTvpUs3WfX+mR4ILuP2HfsDhGfKb1b8HAs+TJ3It1krmv8yW+kynsMMHChHl0hngfbig0/xlFZ6+x4ZrAtBZtCUWCfu
1lsgSBE/OyNOLTwDiH3LVmfk5k1KEqab1CaGBXN/FPA5ZYA2warxaugtFq+Y3YcBR/QNNQEzFRq0KygXgM66VDaIMJi1rSWVB1huJBVPCNaCamWJKjUtbaGnl5es52DN
Mn+jDwctqgZ7tRrgsDaOgAqCBQnROzhKKuNN3TlAbD/dSNooICfj9/HXQTBqSmr/4EoKl2zHQdH2xG2XPma0xJLA9ZRC1R93bZsQ1IZd9So3Zwlk9iEJ2Hfdn8Zlps/x
HzQmN+QFMvNVeR6qlUBSDajcI0STCszP0CXwW2mdmAt7gkZfBcxChSmDUpw8SHvoZdwSTXzAyhYbmbJIsvQpdABRCFOcH9hakclTdTfAmgMOaWAuslDn3fpTGhP1+rmS
U9FX01SIUcBMxtu6crT5JGACZkrwU6J67k9F3lN5BlAFNdf4rwgUaTvVdEItt6x3T+wakTDN9E3WnlULCCSWzselEdEMcz6XX1hZ0fCfjF5MYkXzDOR8C94Iwl0JOF5P
1QU3F3k3+08rgTPskV4wdnENjYKMLkuDsnx53HTP8eXLIMdTObG12BEj4uv+kh3Zr9+AOl1GCRETJl5XF1POMIBRmmuunPwPJ/opox1bE0eOeMIhc81+ukKUgyn0ijFt
ujEkkmFntLtNU3PV1j15S9wZEfmmHWND8DqOUgMqxqF6taM3gjkJG1RVERbxu/uH1Q5KnS76yRkBEJe1ng1IAbAXay5c9yn3uuE1f7IToMzN3HUwDhD6NoKM+14Q6dZU
fsi9i0lc4Wr8jyowUN6FyMCsNhaOZCTfue5oIz0PojDpXFExXPq9IjzVKz2hxrfHjzSk9mlrStiw89f9yuaX8mut4ehArH4ZckJAeTO/OzvKiCbRJr2HgYyrX3ljAm2I
ZJZQI5h7nTNqezy5ilpUsYPwWOS4X4e4usnB2PQWk+/l01KpWfCxArJ+Vyq9dJjN2lXc02CaEC1zfcR7pmqnRsqIJtEmvYeBjKtfeWMCbYhSBzQZzdD29hbUPIbHQRg7
49dt2tZMBQoVGvMf14gX+pkoyhwRG0Mb2YTnq2jNp6O4RY9QjkTlqBZGcymNWvMSN4bbu4FAz8C6dR0hI+/50toDcny5u0aNmVqeXX0LxbLqtA8ECD4B5KMYdQtfuJ65
0F3haYAxI2PI3FUur+Lc5XjrRhseDzFCz+SDjwK4m5dtK3h83CYDArwASmqYHWvoyesHrHUus8PQXrmGw9JzJXQI0bWqh4DiT256h8BWX5SJ1PLsFJPMYVnqWtOW1J+L
EEdLEpSGz34AqivmPJLr8XVhzhHxtPHAQbU2x6fETCzfiHxDz1JvXohvjoz53ICTDar8ZYToAEG4Q1snBUqyWAAfC5CTm5EPA/GhbvDP4fWubKW6aGX64gcUTlTfvh+Y
TLzF7N9T7dSV91r4FsE73pDU5XMhAoQ3hBJLvryLfrKEB89+/w1TbT0H08yeYJbFK7VFI1gz71MFJ3Um1wiIoT7nJ3DkUU1388230SSR9TuyqGFgjmBO2Kfc8ihjWL2V
sWsqCfv+u5Lf4SYhFsq1nRBHSxKUhs9+AKor5jyS6/GTn15PAi8fUrxuhlZr563LF1efTc7asTiV7c/Kkt3caAsj74wSBe2/KftCg1RAfxwyOS3AlxMn+clRctaAq8EH
ZMktE2UkjPsffp1m7xtaQ7/Lo0IEe0yosNRaZNttywivSDYtPh7Z4xGgOSEEuF5jmb5+0wNleV5GuxIPm2/gyejWh4PbGj1HPiGDActwLQgkNHQjBn6P8P3OpKjSyoC5
mgaP2JU5eVQVVpbYwms3vMJp/hn30Z8xcxrZ3IwRtORLLMi1ipPh16rIyqPcGGpSFq+yVFXSFY48P/mIzhAjR2TOfTvf7oxYfi7pNoSeJ6NOn5nf4TEnlnHCjZ6BMVPa
VMmmDALEwjJJekX8+ADt3zI5LcCXEyf5yVFy1oCrwQdkyS0TZSSM+x9+nWbvG1pD0F3haYAxI2PI3FUur+Lc5V9Ty227SM43VC80dWeECU0tfTN5aLqs4f/9pPSdrJHJ
lwT/0a2hUAfsP1nJhPU5cfOD2K+JuP9s+xpugOCCL5Z30fLQlZH8U0qd0o3+hFD3cmrxseG9+jlp28DbjI/vHYgQqiWa6qIJHH0RJSQVQBm29TcqMI5FOpZbPfMRnJp7
f+CEcT80jdXgbbECTzioeosIP6aRfuU1PrJXDiVxIOVwNT2Mmrqdmy4lA4Nglvm9BuoKHZ2kYdjLueqqxM6WOoUm1Hych9dzdvsM36MMB5QpkU6xFP+OrkzJhGwz4IFx
jRHMM/c1TWfwBovbUWZxCFaiQizjjoois8EUTuBDO0x+MhxtkNz/FR7uCbwm736vN4bbu4FAz8C6dR0hI+/50toDcny5u0aNmVqeXX0LxbKTfSeZAqVgG8iFKlrC8bHe
WHpZTWwke/q/7Jb8J6xKyX/ghHE/NI3V4G2xAk84qHopDbeq5eFsqnFW9BP40WqF1Uu5andBiNIrgpTZrd/o/We0kErWVZYk9M9hTi4H3ExNdBsVec0vO/aD66akjta7
bPgyCvKIXnStbcNnQ5KEfxBHSxKUhs9+AKor5jyS6/HIh4yhKP+L2Uim+QUsB3CW6QvkJZ5+nXWHc6Mc/6lwiOrpBKzO/Bf3KSdB5LIsN2per4RXLLvh77lNdvj+IGfc
uOPcwjOEUgqSu0W2PUkbuBZCKEf0Y421uj+N+ihvvBeo5xNuwlxysDz/TpW9IRpuYvE+ZzrVTIWM8TE4Y43W4YYSBkyAVpqi9nR9Jx9OTIRKBAJIYQG8P3javccq9CN2
P5cEM0RFQCu3YUfFOGYOCcCxSHencC8/dNmWzL3KMJj1b9G1E3K4cBsp8zBkeHW/JEx71mMBN8jmcxFZyofjQP/pPqSf9oCqNYCnZk1m0MtVr/ClIS8L8ZiO5mhu0ceG
yesHrHUus8PQXrmGw9JzJXQI0bWqh4DiT256h8BWX5SAt/flJuLfZfsx2aE/2+G+YMsXZ26/BtP07qChQQ+ulJY6xqlAKsRbGAyfny4BSMdlUJjKIh86lIbEuBo5Q4JN
Lsi5UI13ay8RBCw494OZRo+ZPzJfRmenKzy94wxUV1L8CvFL9nXrqXZvAioIb0/7SEJclXkkzEA79DYQGfEZuN+HqSVLw+oyrJ+tkf7N0GVndxIa1woB5QA1olE4Z9qY
sIcvvNE2xczKiuxEV0yFjfVLGukP9KkztYVTHggzD9zVGjPxlVXCc33K0ucmU24ibPK8EE+tbhcKjFzl040pfHOMIhigMjejTF+xOskhOiT5XIyWwuGOoDY44YVj5r9K
pmUhHOdK1J9LF0HBwg7Zsj4j7g1puFvFBHCWHh7Nxi9zK5dmRFHjUTsk3By1CcQbU3eDSGdk1YaxBG7QKmDCiwAkLEg7gm+OB3+rjFbTNgCnnV67NawwQGo5hfMaP2T7
ihczWMAEFbOlWqxRb3+DM/pcAhCm4m/Wsoxb68X0yg3E0A4Yj8qtLZAbSzfO2lGK9JMA8cgSzw5b+CVj0ranGOXmMphu/1EO4NeMuMgDrGWBSe9VGsW9g5Bgf2y8s6U1
Fz6ouR6IbzRRSydezSyznFQCzjR41ya7Y4LPhs2BvSFmwB2Rc8N0XkgZL2LRlejF5Vk71UGX2LpxAQa2c8TcjyXOpG403N+S5xdGGwMGCuVZhxk1+ja4tXRP9hR+kmBL
hVM+OJL1tcZpV9mvzYo/dQGyMNJlyhAje8WxUJTUODmBARWMAL0pWixQNZrBij15cUwspjv167qSzQOMhncQYsnrB6x1LrPD0F65hsPScyV0CNG1qoeA4k9ueofAVl+U
5EAT1KzW5jnAUJoICH4x27vtT03EHCTxSDAa9NERV80tfTN5aLqs4f/9pPSdrJHJv3/VtFCaXpINCeMPgRIvwUqE//An+VukiifW2h8ZGg2JCuyBdiTbo6RoMrtgCJmZ
/3vQwyp8Mit6vANbO1OFpmbAHZFzw3ReSBkvYtGV6MU2N2e5el+vU6VYuxGAixPqHpgJCrvZm3662rv9mvTCnaIBBgNdVbxIaOLkD9pE0F3AsUh3p3AvP3TZlsy9yjCY
HMnE0W+7WRFEXL8s/T4mu8ZPOWrksOQV47pUt4z6sGsp5WZoEFFrlU+wsEpR3+m6vhc1OJZ9B28q4Frmu73ZdfpBKXxHZF4CuX63IokB7D+C5ZwP5vMo3HEzc4WFYOHc
RYhYXhPQS99ZfTSaIk67q2e0kErWVZYk9M9hTi4H3ExNdBsVec0vO/aD66akjta7eM9/W2mzzWP/vVaeCVrptaDZUAVW6csq9L8xR1CBHtrVknuokoPXXs10wyccBszJ
Y81TpW16ZEEBpCit+g7PITh4Kssrm+IaJNjFJVdCFVkfyd9yVuBDtqMKuyEpvdai/ArxS/Z166l2bwIqCG9P+0hCXJV5JMxAO/Q2EBnxGbjkRBY0ru4IHi8T9ivzM1GU
Y4ChjS2s1ZiX8iB3fbh4CCnlZmgQUWuVT7CwSlHf6braNbUWZPBSp5VGZ89VDmJqPfigjpPAQ0y5qlqmsDLEQ2U2+njo7lfm4EPILSrDcLLFGM++50nwJBizeb3lXj6E
Bbszhi51AbyQxQoWVVEHgkpNX9WO9YoDwYg4CzqYrMvs7MqFAO8fuFNYu/OC88JcR0JlEHzX3CZY9syZgHzTdl2wnlmOiVIwYggkI4iCRgi7uunaGWK8JajlzSUtSujX
NzhD+5IjBRz0vETmQUiF3mHZQ6EgaTQPST+v1NFXZ9JpS8zC6MLwecMOObdQV4lZ/3vQwyp8Mit6vANbO1OFpq2dM4Daxdra71kSImyPy8HpixTNk3nVmKEpE4LJfmi+
T6bgmUhsGkevbnpRJgupZOjYgmR6+iWsEb4lpBfebTbWQP8KF1xDuCdEW1vSWkNWleVPNUjRjTevattsgazRCDpcrU2R2ToOmmXXCCI1SK9Vi7DXpwNsPeFw8RO98j89
XPOyDk3IC0mk6GbfpWB41AgI9Rth/wlM8uCDK/EH/kERbnd/CRFKG8XtWcprYgASkEloT/cWdx77jUQ8clNIrlTJpgwCxMIySXpF/PgA7d9ycPFY9ogtOHx8z/sVKJvp
YtlXxGiLkGka6f9HtTYphAOJEb52+yMDPSX/2KgucVR13XN6EsNK2RH6eD71jR5v00TCo1N0I0pg4bMAyetptlkc+KluFshx0AQbYwAMfOlTRqua7Qe3uWp9cBGWcZjk
ZPqDSeoo29r6a0fDzjsiLe3QFm6xsylkLBsIfHb4rHi0Y8HK7Vw17Vg4tr1g2921yogm0Sa9h4GMq195YwJtiNNEwqNTdCNKYOGzAMnrabZyzhknjJ/uBlY7U1i2OuqB
VDRX0pZbRYSaizBmAEJ1DZuRfpYiSIxZd7pO5V+PztkcwIq98yLaw+bYUksRkofvE01cDWsazdnJMv3Gbx1V4Bsj2+SUvSb4AXXAWlIOLVJYellNbCR7+r/slvwnrErJ
zKcOOt/zGyXVZDGVnzPUpxAwMBCKx5OiWVU2s4a4IkN8PzuQBDSBIpZStjvRXfNkStTSmNes/dPNs6oTxYTaM19w9TtnVvfoCb/mVWJiWt1gMcjtaSQ3b6gvvk62lSra
mCnWY0weDJSNyZzPWqjC096iQVfHG30+H28jMPYp2Us2gj2064rnD545hdtKwfgidgd3lDBzw/S9t23s6niltNBGBvIShjWbb6xM9eJ4upb3WrIuKnQwnIhG4gUgM/C6
adJse3ESmdIDZN2HCR4DMfdasi4qdDCciEbiBSAz8Lqt358n4naGUbsXTfxUz0IlVVdF4dRdtkJob0Zw05WXCeeQLxayVInjzVH7X6vOxlCMvceyKd/BING026yOW71G
nANjmG+vlWLQS2py54C4y4NGIuWXDZGUonciZjbhkzLza1DcbhVLQKZvtb0rqqPSBATrnbW6pUaORi1sTHdPK/iA0DRj7GANeqZPCVT5EQTZxTYUuBX9tfm1KALH/oEZ
wk4GjEg9SmALkkbIFRyLmEt/BBIlTo+GemH/lE69jShKVlFmFlZOHXxPDTvy+7hWEFn/chRLEU0wyFxhC8QSg5C7yS90NgRAgGp5SgsSERaDRiLllw2RlKJ3ImY24ZMy
CSXRgKc0Zb4JKBjhONNNsMAEn6iCRzS4G3tdBwIq4wVHvRC/LPMqlFDmLTb9DFOVU0armu0Ht7lqfXARlnGY5DOWVJfpO355Cs8VsDynAuoWr7JUVdIVjjw/+YjOECNH
fb0nE02kX+een/kRbqH8Ju93MN4NJdo3nLlbtMFvWDsJXcT6PTzNXoSNQpwCo/m7CGEvIQKFCreEdBVaI6oVmyPu/7cgyzkOwLBljAowRsQ2enWKJVIkwvLxd1xVt5YV
VlqTe+kRZvAIZzaWsnzQ62gRnu1mqPEC8NWYKyTyQ26MPXkk7KVBQqcO050UxAlTZIeuNiqyZTkOsY+XsHmEMjHZfJlrYbmWT+aETjING7KfqRSORCxjDx2L4pyEaFRa
mR1j6wSoabEG3IBIEMw0X9SQh7nW0KjLfYpFwPyalhpx9PJincJwdaxM4emNNZnFKm8L5GhgH8OofZAesMVw6Pn+Dc26csCzyEFQrBZ5syv/XUswnGAsOyDoD9J3sVuX
1jWCMcOhZN3qA8FObOI2E2fP6PNwSfeLN/Xdbi7D5i2cI/AZvOPyScyVdpDxxHwA1JCHudbQqMt9ikXA/JqWGjiuzYrpYApmoJZezc1+W+cjZUpY4/x+Gy3fZeS4jums
GZiHVmm8lujwJ76nUbYoRTdsu9sfVPscy7hG04fisL2jkxWzB0rym93fBkp124ZhuZclCgwQOO4caCs8fNTLGfUSDvBLS0yBYW/M0cA4K0EWRKLax9CrI0v9rBaRkXoF
8ZLI58EBshuPCqz+j/xjxBoEClaQOE8mYmklAVQvFkHEOG8vLbzdviE1KbyWmfETvjqOZ+f6LdSREpusG8L23Bx/jsrswLJN8mYdN5X2030AdtKOOVodm+5cyUMq5NpP
CoPJxv2muZ5z15OriTJq6BdVqlJlBTzzEA/Yv2HHINTm25eNGN2vbOBzRw5sU8IGaMud7iJ+MyoRtXsJgnjalnwlPVr1vuXQMglexD0keNv930E9P9eYr3RLruL/opcm
SK3HBBw81b4Ow0QBslfAZrjp+Pxazclc+lWuzot+bXdIcO/ocOwsHEhzaFyR3c8ATUe1826QekQ63Kh1PV1bIhug+fYBaoY4VVxsNS5wssz8ReAjK0E3kd9UYcj4av5p
gULEsM0+JpTKZBaYo5fsT7+n0aOgZDO1d+DKWe2Ny5XDsYqM/8a0W/Frvt0ezilSSZXdRwN4saED/s81w/rdTFmzpa6j8B/JTLdjyRCpnKoeQqZtGemjHIuYDigb9rfE
NWF7DyP63+J8sQLB3ENRHkitxwQcPNW+DsNEAbJXwGZ2adgKXLBEY87ESGg/aLCOJNdJQ17RJ/R+GwqHSQjQ6frDQwSm3oe+0dswzT865UsZKIyrzcDX5xzOosO1igOv
mABiqHJPeenQv2YxmUEDz3EB6+LpmpOMFagkLUaWeGkKggUJ0Ts4SirjTd05QGw/HVBnWIFtnkdCLBkFFglHx6EJvxNKzAR+q2vlw2G4o3NOUwgccYxhN4PgsiP5+rEw
nVxA2DCCtygSM7SzZu0TUhndHwZ4Kaz8h2NyrjbG+5g4fp9sZwofx8SO7NTogVX+JUko3yFINxYpKdeSPDVFC+IF7KvEDlMteSa6DO1pae5VGRWnbyVf+ZfwiIsuZl/O
jdevm+9RQutkYafhcn3JZqxyJtlS+3cBhrOeOdAkQDRuyFV1vlJKb7NQSLBX8CAiW00IASHW+4NhmkyHTpCGUUitxwQcPNW+DsNEAbJXwGYLn2X4EMGYntDQYnUosbAz
a6NThYSRL4JudiHAeVeXLtlHnQcsRHnvqwsl9PSAtIJsdYBDWAV0rU4WKHww1KIinq/EUgl9lUucT/rS+Uk7VUdwJ+7qRu4BeClMc+Kacvt3OVvauLBH+dE3wOKf/ERG
i6Si5YGte2ocyn+fjyAT8Wx1gENYBXStThYofDDUoiKer8RSCX2VS5xP+tL5STtV3pBFMW9m+8/IrRoTUL+WH9KdwBb3sv+PzRWz15yRvGpsdYBDWAV0rU4WKHww1KIi
/A5XALi69MADeB9iZGVgHLhNIqH/m7U6kOS2MUh/CzH8qGo2xYU4E/fJ+5uuWcXoyogm0Sa9h4GMq195YwJtiFzPxsg43xdL7l1deClvP9xVSsK0WmEE8RWiJP2HNaOd
GDeBHnjDwTc3ErFmpNJnBQDC5atoe7qSpzKLaVXolagM98rSoDrOqshq4dBO44rzjg+3U7w3n6PWcX0Exy8Z5shPhxmI5gZqLA9gRoRY94/7oZsKbDqwCNYoiW/zRBgI
`pragma protect end_protected
