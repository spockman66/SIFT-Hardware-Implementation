// Copyright (C) 2021, Andes Technology Corp. Confidential Proprietary

`include "hme_uart_config.vh"
`include "hme_uart_const.vh"


module hme_uart_top (
`ifdef HMEUART_UCLK_PCLK_SAME
`else
	  uclk,
	  urstn,
`endif
	  dma_rx_ack,
	  dma_tx_ack,
	  paddr,
	  pclk,
	  penable,
	  presetn,
	  psel,
	  pwdata,
	  pwrite,
	  uart_ctsn,
	  uart_dcdn,
	  uart_dsrn,
	  uart_rin,
	  uart_sin,
	  dma_rx_req,
	  dma_tx_req,
	  prdata,
	  uart_dtrn,
	  uart_intr,
	  uart_out1n,
	  uart_out2n,
	  uart_rtsn,
	  uart_sout
);
`pragma protect begin_protected
`pragma protect version=4
`pragma protect vendor="Hercules Microelectronics"
`pragma protect email="supports@hercules-micro.com"
`pragma protect data_method="AES128-CBC"
`pragma protect data_encode="Base64"
`pragma protect key_method="RSA"
`pragma protect key_encode="Base64"
`pragma protect data_line_size=96
`pragma protect key_block
taRoeU6EL1nGpMu9irppXN2mbm+l8MvKBEN9TE1iYB3+7+zAjOG4gtmhjGqiTj2Tb311hVPSEtcdEhV3LKF/4KxseSNiyjHZ4lOyZtA7MQCy/uZguJ4s7g/XczykfMEV8icKbaRnxfsoSAbTuaR7ILOcAd9JEDSVnKONZeXUFCs=
`pragma protect data_block
IPsOtGCwpgkYjw6YVR804HQ3JZWImrB2Lo8fOpASQMsZoapVagyXVYaySGYzwXxcQn07R7l7eKoSKOSpbbYZrB0PO8KM1PvuLY2mOQA86bx8PUFsEfxY0pKu9/INpytN
a45AQE+CvRbtELf1zPnpohv28tskmL0PadbGFKGK1UsdDzvCjNT77i2NpjkAPOm8DyRwX8zhkVFTxBRQafZh+sTNU9Pbxd20omFCncRRTvduFBBvs2HMdAu/G7k22ifk
lBoDJbslkZe2it/XYpFqBzs+FcowHIPWZY/nMBcBQ15cTWPCN7v/RdBeQGPMqjygCcrbxEQRrfsmnDsAVGjpFzu9As58ucoYRRq60QDPcpj9+A48tkgLr/QxUVjyJWAN
88Ql1uKbqZky6rAZdX64cGkVLOgeB6P0JF5cx//ISIm+fiq5YSfLKpI7peM5WPXok2mWRN10vGC/4GEmsk0KePsGzWnZwoL3xAa7QebnSpegLZH3fNXkAmvbvUOzLtpf
iRyJ1jpW6/baJ5HJNgWuyI4qq+pQPw7Blmc8JOh5sXlMgYvOqlQDiKKxRZYUO2XN2RSRGFSm7XHFhiZdlmAk7WqL5eupP6OxgrxXbderBk8dDzvCjNT77i2NpjkAPOm8
NsD9+oM0ibDuMFQXYHpe2QxiniZr5H2XUJZIaWWWxx5LCbH84zdgTjfdRW6D9zCiOJHO2Bdr4/0Yl68HdRJiwDauEulE3MGi7vZAivr3/BMSnUHMIUXTu71O3cC5kQGp
X85o8TXdE5hMUfsa7FyTdu9Jz1Phh103cALffp/PlHx9Fqns3GzCzmPwxl1E9oZfPiIf2BvOih+OWTFfp7+W9jkJ/s9u7Gk7H+f7wRicrMZrMNOH8qbmfyEgz6C5HzJO
lSXZ8lPw63vBEw3Zv4b/mzU1aLSAYEXZENcWeNxZn1FrjkBAT4K9Fu0Qt/XM+emioEkDTihuf52rvcOZkDX3Q2tqVd2aCMUbHVkG2iWq6w0Sp9Suf9SKlhlvhr4z3GWP
xJIGQlTD/zrtxY3bicvJTAN8ZKspsuBlEc6kogTD/HJmmk9hcobVGxBWqFiXrVKSkN1PatxQLn6ARD8GGEf79eCGlWmOYV6mqUfKc5fG86UXGLQptCZK6ouUjx04O10r
1vvvh7U+VOIjGctapibyY0dsTxHSMe8UaREA9s/I8YFM7U1mvJcn7VgJFB7BnpD/rZY+XdSkH4lY6omSSWNTVxSH7XIL2xQDZyHqDAgyzZeft5ZDSYRfkdGMXkojQsbL
MusH4G7ykXCw9dTlqvNq2HFfVbSXc/HVQyHLgwggSNIOHVQvuvP9ruTnzXEnniM6cdVxAOf7l+OfRC4dEgia/pDdT2rcUC5+gEQ/BhhH+/Xb+TzAD+I++q55UdOWPD/w
qg7w03osV3q3/l2i+eboiC85SqOfz+Buj9n2HaMbdFmZD35YhCP6MBDUBQaVFeInA/3Juu9lD7VYgD606D4na1iCAMTCTkNYPMHHDtW1EXszCLJCcjmsZmjtO/0NhZvl
V519EGO8joQmN2AepdazcwZLth4sedTVe2u9FXEDvDXwLaqB+S3orrCAzi1s83MqajmE1mTMfqjAr1BPjhIDDVs6/C2A5OYlE45eSVm0TgRA3Twb6A5BS0jhmpqTWoW6
DLVkqHmPcIexgqfw7mbLmkdsTxHSMe8UaREA9s/I8YGLwoItLogypANUrDsB2Wl81nFKXUBKNowlO3std3rcdqNJRnCwxiTvfu339lbtythHvHh1DmhfixiP9ma2TDZR
8uO8w9B25JLsN7jRqVQCewJR6hY5txDXcELMeuwdja/9dWzKA+DjBeI3dp0eRKA3I+hcKmHH5f4awWtHaJkI2PROhBQfpMTPN3iVb//n7t8dNbZ5fXtLzhbTcGq+C6Em
h+hkmzBZjOlWNdS0i6bLPvmRO/jVJmyoUKWnccN8zmnqmd7JXQ/A2fQ/Ev0xX2P7KkHTYLZ3eFVgR6Fcq8b8rKo8pujVUPbagKffu/VWf7VDsZk+DNq4NWo9oXXS1Kmz
9jTZGKJGaIbRJOcjj0vuyZDdT2rcUC5+gEQ/BhhH+/UUwmTY5A0ncwzmB7rB6TZBwnhpVTvwwoJr/ftGExDiE94F73gb9oQZhAwrLrz7NXEQ0YSM4fYTWCRcQPGbx745
mVADzemKIvfhjPmP7tT2Dnj+oRQhh8rMQ3EVD5iny/cqQdNgtnd4VWBHoVyrxvysMt0OwKcA9Mto4wQ4LptJfvxUHvS748xbBic8fD18R50cyeU44S+8TsauCKwl7Fbe
d55E1Q3T/wSt+288zGULCmRUmqRfecW4prbjoBiJy95A8V0go/dR9FvzMBOO+nx+9gU1emMfdOh58qCTq8T9xZDdT2rcUC5+gEQ/BhhH+/Xzxf6mlP2CP+gdw+v7sNbq
UoaSB4PwCKWe1YVCe4ZMN/2BYN4L5Jv6vF6dovXyqr96kMFBjgO9EZXrc0pZNwIiE0zOG8Mns5Els4ALrw9FAq7IJwfc0o2Lng6NZiBdODl3TIy1pWvpGAqbHdmoSzCs
jIJz1JGHnBL/2glpQEv5zskQHmjlHOHeq4CPcXaSZ7H98/imnfcBjeAv/NVwupngW3qoFY5nENev9TqZj9MrizHK0ZM8VhHM8+JFRIH2iBOaPQFQnPm3H2WDUYZqTBHz
oZ0R39Rao0L/MQGa031XXErCzuvHjgg2Y3qC/PxX9ivJbvGdpVDTe6lMgc0nrBgfkGCDG4PAdUHCmYI2WUXquKdykisRdBh98wZaW8s3OveFdO85+y7J6sCEnMK1g5h9
Sxzncq0UE0mV1YkTTY3dasutxbcCIbHHQqjzcpwRSY7CeGlVO/DCgmv9+0YTEOITG4qNXrXEwFzl5BPt30lSLEdsTxHSMe8UaREA9s/I8YEfdT5zJkp9QVQBPEZnq2FY
fWrvKWjV5pyYWDayQ1U3k76VafigQlq3QOMxrNep8jB+Hxp7XnCfIGjyWRwgdkPqvpVp+KBCWrdA4zGs16nyMAEja0NrQS9enK/D5dYMOHKoEOb8/qjEV7sMTEQX9cpS
vW5EnQ0MG+f4cSPyLjmGCEdsTxHSMe8UaREA9s/I8YGHq9ib08dc7Bw485mhMle0BZMA/e+oK21G8fyhNo/WzD+nOccSSria2WgxULFY9SJh4YAPvw4jNAzwO9MVn5FF
vHcinE8bUQGVTOi3NIh0rGlDX/EwREU4/IdrggfvfOeCYMtgWq2heSMXTXF4wFXFKkHTYLZ3eFVgR6Fcq8b8rNVVAhzph/W3Q83++xOW0KhPDA7oub98bVjvgG+0+nMP
NOqGqg2pN3+VQcgXp4ZJWMy8RWTJW7KiisSsD6uE/F7OMpSjdEzBme1bwHtcDpcvBzbc7D9Kj3ZWu/WOAWe+0Ge499TfudLj2bZdAvQ7ZaryjCBdRLjBdYJFUAXfWiZD
zAfvXGnYjp5E0NJU6HLxepMI5fjTTWWjdxoFBzTCPFre2DfolkiNM3wPtVD1H9Wyy7IGKClmFz2zNoK7Kymdpt7YN+iWSI0zfA+1UPUf1bIvd4+AsF7VXN0OVt4fhbwX
2/l/GWDGdlcQIVbLlSMHXv42kh7ZXzlHS0s76fOTvZoqQdNgtnd4VWBHoVyrxvys6i+ShMstNgVeTreEc1l9/AVx61uzqPyd4UU+rJ1kfTQUbdvyy074oHrSybZzPI6K
I96FziJ1TFPJgt7N0D0zp5YE7pGr9oIn6fhlX0HZ9daC1E7QlDUUgdF4y+eMy2Vq6GOujYR6jCcpStFbYTQslpEL/qfj0I0vw7fAsIGmcPXe2DfolkiNM3wPtVD1H9Wy
ph3G/Qj+f1Pw4NiQjkyvY8J4aVU78MKCa/37RhMQ4hOJv7yiOfD3gG0mYjj7Ngaq/FQe9LvjzFsGJzx8PXxHnZM63NnwJFbl+LgXY89HrNd/kLMk0hyGVBPsN6HEt5kA
v3YPoM/fU1NgraYKtrkpoNVTNw0Hz3geeXRCQALVWp0KTqUGCcvqA4Mjs+te4NhwfqZV5yGSmhtEwb+d6oLQYaVJsOlmftgvDRB2azpqXtoIVE08Qtg3g2g/g2Nwzk/S
JWp9XckB5OsqQjFlUBkBYfravKb+LztG4UPfSILgt2mEdd/Ur3pqxnHwdxOIanccGZoyC9WJT4UYwh1M/1l/klEmb/PljqMgLmrG//LpA9XA5vBdiOI7Wu/3mG/hvCDR
DqfKTG2vDDyPF067um7LDk66IlT/V3h3IGLXwvwEbjEjDXdqy7ciMmYC+dnTnjXfLFXrZdl1ivE/2ReBSr9N163gYkcw/C+EyZsCfn6cCsrfuPZhesAt+mRaLGCM7JQn
M6/Lre9ZFh45LXqRRPycbm9a5o8x5/3ndRZpvWL4Z8P0NnhbOwwnl/wUBWb37Qn3SUNzdiTAH8bcYYwsp7tUSM25QN86rV/RJrtri6oSPQD5uaDXgOSnEjq2efWYNte3
/ppbkeDR8N34ZFPcQUaY+VoMN2g1/YQGanRQuK94vApYLHFIY1RMOzlk3TTarlQo/yeAf8vpnl28wLLrqkmqzjkDip+kZoHGAKjICF7nlCx5iHKQJBYRazsFHAslmHos
hdjNLKBApICFdMzPCrh7N02s57Q86Wae8QfMbcO4Bz62hQUCRuR/XfCCxrnAF4r45UnMcQ2VABcFsZdlVhwo6Pzivb87+DvEOYlqgVxEXU4xTfikH1vjNDMuv7emSqQf
3+nZzd/JHZ/VASsMX7plupQs2bNh8CGRwj6wiEDW9q7EvRJ7zeoKQW0BCD+XxWsGBcNy0xL5JpHhqyY1MhBRz8EzXqWTpoBE78SFPVHAZJ07LX1zd4LgKENs17aIZzlz
s4hMCulksXCNXhETnbaBk4J8UM8ydLRwzjsMMIVoOHzxm30fPLIgKdDaKOWZg9790bnq2cNPGJdxztHr1hLFX04eS1kG2APd03W+wBKqxMh6FwJUrVksp9veRs5Yi+j1
xE5CXlC0wNW0El8WGuPfjtqm5rD9zAkgmIvDD3m/AgVkUcpvf0uQKtURdGmuE564KO/RnvaiU/j245cBfT7ILVW4ybTErWMuWtx28A/jEew5VuM7PKYP8oXMQpGSxUH4
O7ICGC9Lt0UsPAIAo5ZIxv42kh7ZXzlHS0s76fOTvZrHWebdlND4kHqJ0mURTDEnX9/LrsORNG7lFcJ7o1PBowc+FFTIwjeHq70DQTcuIqEzfl/eN1II3q+/jCQueSIo
+nH6WAFh3OppoH2WP2YIJcKOZ9t6l5dVjGKrqaqxdOLpq57bVFPn5gh8VmCi20tgWG4bTxSnwLTwt3zL5vHZ3sNJ5mPkof15V58Ag9xm7feVdGf10MOfChw88jZq4IeD
d2Rm0AhD2+a/p4j1qpPSt/r3K9E8plDtZ0GOkGEy1FK1tpGvZOqkl2PDAIqFcBDXxRKHf4Sfd8kA7MrQ1CwkEoqrAPRVgAdYIiPxcOEeetVz+cPMJyRaI91t5RJa+6yY
5pQxck5ZjaOTQiOfWoYAvFa0rNcRJ0faCB+q21n9n/csQsXKDx4kauFWc/K05EH9HFkSGJVR7qls7wWZke8W/qNVl9IE25jd7tWSLzuoxY9jU2iUtL6D0teMNvRDvk51
1cAQhMmOga9JFMX2gqvBFB4hPd6+4dy9I0YPDQAjhwcMNJY2Q4513weP+uZvZl7C9r+tL568IA38eLxTEaQpvgM3k073GSLEUEezNrLbAFf8Q2I7xFiVMoWouZjudZpQ
BEBnJmy99AlZfuGJjjPGQjGeE4qypHDDPfomtLjKfsb6XtkmivYq8EAZ/kDKkZrUd4DnLVka83gnQwSl4Q5v/UzDvwDYX1VwTdrNEBAYxj0yZ+WZLW9GKnuXv3cXqsnh
n5IlqzU0IcI+C3Mva8L88FQR6K8Qd+8w/1wORAmI2FP83Bfhn0WQ8/9L1k+UBFNEQp/KAQ99DyxFqyH+oJRcaiv7vAIclxjjCdXzc7balykCOC1cUb7f+EwzpJ/keSzX
6lTLr6sMO/9MBD3WE9qmjOdTB+l4XjW1Aoe4kn7G8ih8q4f0NbJSv2q02Q2gh4VhufAwMZwqgomXJH2Iy+q4pPBJwQE17sbPj/vPIBudbInar8QiosG2Tcr6WZMLF2g1
LKh+WJPBcBnxQNF0xYsGuhdtDqj7AEIp2VN+QzOmBWXXqXvDgV/y/A97WkbxMN14Q7JLZrx3Fj4XhsOxdJeZPhIRdL4ItNHTL24qhgJLs8wqvw/eEFSRtHf+BmQZ2Ppl
F20OqPsAQinZU35DM6YFZRnIyJv0LBvTV9fdDn2cUs8racBlDoc4P8n93ghyZ6qJKufaC8z64atPOMRYN0cfJ+bSQ0jl8Hv+Lv2RIb8fPw2IKYw5VO7PNAPBzZ1KBfS6
h7BY3zNCKMOR25LsF9Lysucpckhr4WKrKVI4tctHd2HluI7PrQ7BT2y/sAf+cQkdpnXQURMiTn+3KF2B3VQzkYgpjDlU7s80A8HNnUoF9LrEik11wjIwlVxBR/Y0YcJc
ZJ43QF3kD1wIDY8Ts3QuX47UzDreiuyMngQmqyEzJgFj386pSJ8jYi/KOUvPuTVLBwgOxNH418nO7pE2b+MekQAjQtFcwoiwTGa7+Sl3Egk1+RW+kY9skfkyCA7oqjuW
FQ6Z/KCevA5CWhpnzF1XuM5Lf2oebksAl3Y8FKjJzUiXP3xB79ycAR545nE72jSk+aG9jNZSQfIivhXVsqAJIRBkWqm7mf56trI6PeI+OSTDbmeC8R1cKNuYtbZmYmQ0
ZahePBXaTrpqrJBnKOweIT6EX5aXQoNUWnlW8ddqhkLMR/P2Qb6FVnOaoc8ZT0JlAvxGVp45f9X3WFliQvPCqz+ZzWmcmT/LTSBvMVRTJb5aj5yakJcrVpcZ/K5jN00o
CPmSQc4DQeRK4oXOdgcGyobno0fCQqhgJ37U+ZlHMW5HfUsOXQeY6LBRS2LTf4+Oc+jKxnf+qaq86wXLcHjkNSCqCB7JCv8kB3Vju2JLkk06noQnmD6wjzntFcztc1OG
nR/UrlYayiJzfcZOTpsSTpT/nFmox00oR4WHsZyNw1fpw4aGaSIv5dx7b4rUsMFkBrQiJfll9txu+ob+M2wn95OSGvbwSgRQ4C/BRlmAZOwhON2sEjjvXM3ifhCLMEA6
U88ygT4kL5EpOZKGeAPz1sAF6wo6g5NbDtOmxImMtoUf3ZxAbT6YJW/LGPeHDekqVvfbMROq6sixSIUlGrPD9epZ3HQ63ytekuCJffQX9jf//QgdZMlc5aJ+C8KzMUij
4scqAs/SZudVDhjvt3JQywG8en4TnJVar5jIPXACRerh6eBUStSb61Jkd5n5nZUuRTaD/GUsWSUq2WespVEXRq9aEjbomeKAEONBdyYGwSYGHSeyiRNS68ISK1gIGybE
sgxSHdM8hDWr5RvC1u7478ORID/2Lv8NZCOTiN0hhfqTZC28zSYilGen5B/qvO8leffLiD7Ac3CaVxIE1eqHJbdW8TWBYeH+bXQ2NGN+8tB8FWWl5gzSstehJWBR3RTi
KyXVq65ZOeIGys3+EEtr5Uck8qHr3zrIp3bShAfDGFuRj8PhjcStZGaAFQn6pHhPckKMrnzt7xGbdo2drSXcasVRfc3wz+hZ8iB7iAPu50Q3G3ESRRRpvGrN2dt2IJqj
ztCbrR+TYcdHCh4Owkk+W+sZVf6oqTJ2TyPjHLuvmbrH0mMjDYyscSQyCOIwXo6w16BIKnsV98ADH0HRF1PD58GlZuNY/PKePv76lEmiyh3WuiozITBaV3FE09O3b3gm
n9onX8CIjYRiXNgwosFsJzm5OA/n9lhImebMSD9A7iiMcvIqzxT4OMyMWoa0cZEzuu6vbrhyr5/KFTFzwBOBejg7ZA9cKOCY/9MRUKSUD9qcE3AkTCzr0XJPVd6nUb+0
H7QrcYXpbus9aTB2/kFutdoRiOSq/G3/Ik3qGe1hF2DZ5F1mcpg+SdWLpOPtCsjRBEcGsRovben+XzH4cBVaquPs7b+2OBFY1FGQd+NWDd3S/k4GQ/XJw4smoTtFjQEh
VT6Hc+flTtdd6dKYCbPi6ndhhqCcnmtxUyW1LEjJCD3Wj4/jRyZQIVlgoKXYvSrWZSvmx+Mg2iy9GfMFUeq2vHddwT/zAN8qjrgEEsCZxWppvD0kXqb49sad1dvxZ8QQ
JgYYwL+vZE73oLVVlNCIIBoPhdV8cx9OAvNY1EdYQp1vc7zqXR2DiGergc1CXLrFmf6hij5Y997d48X2YmRGJWsB+mQnnJN+9QKkUrs7ec4yXyOXCHIHIGBNCF4wgnkG
j6aLJIfn0iF1H8ExvrHhEA0KVEMtCkABXa9grzDZQ780LltWzsc8B3bBtzN1FlncjDKFHnqGXX5ruPi0H76Kq5RoxClmgo8Q7OFhfkdyBRXn3L+8GwID39C8HMAW65nh
G3ys7ImtYEVUssI1WGNSbvWNfowbLrinMcz/vYgCL/T7NyThRAmUbsTA4b/nfQFQENgbpnG6qeZ/N0PeS3KYA3eivmml8T0LAFUQS6huHcgq9ZyB7F1OgyLoxPgU+L4j
z4z+i+byIjI1n232vvlz0To1SUZRgSvESVBbMfuOtBdKhDk2Ci6Iw0vOqmPhCFD96xl6A8mlZgJloJFevbie2zhRhNvNgjJ0OyAMqOa+ts3d3nf1y390rYK19blxwSl/
nNlBQs25VIMYOPIYLwxhzeVJzHENlQAXBbGXZVYcKOjIayU6Jv2pAfOU35NoWwmYUS1IKLWX86Epz71VhNBFXmvGQk2tkpNIgAaCE+hKuIaSNpleoP55fR4omjpLtDpS
hcrGMn8593XaIKmkNg3/BWCOxY7LTFCdSLFAzlc7r0J2m50eo7ZmeJiHFRc/gfsMVqF0WrN14w3t2SbPZAHfpHZshAbSu02L2ZvVn/KqlgP5HA86i9SF2A43V8E48lOd
1cKrWSRVfegMjWkdO9cTq+W5npr003cy2YSL2Is2uEPgZiFhMiVuOqOyEr2InuNXVbqznH//u7cm1aT9srGwAaH5VxNIYlmgrjSU55eLQhQKTqUGCcvqA4Mjs+te4Nhw
aNV2ZYBJ9W+lBKP/1w9uWLT1CfcvCd/in7YKAfSoMuUdth+UqoKODo62Pv/tfKnxsQnQJYjSaD0pIqxKNbTaFC7KnaS7rx8S3GnLI4RpW/DVthkC/ebjhf44bYDelN7d
Hx0zKkO6FH7HZ674bNg9NFGsJJkZ/sZn4P09203Qa6/rfJIOBCQYW3JlVVDYsS0UDqfKTG2vDDyPF067um7LDoW8eXDoHZl58XjYj9Ti2cblkCvulf9z3izz8v/oQDiN
7HY7Tcai1bwcSt9EP5zyuBMqBSAjiEf1i7isjPwv0hIIoGKVe+iwVmxtOZy5elzLQje4Y73s+ByuYal9Tf+8HSPiHcLkM8VAeAdEtQgiMKGeEc+fVr/+w0SaX+rluPRf
2gJvN8DL0sCJaPjZsbUyoa2iLHqq/uHQtUcNnsXUMjkyf+1zg4haWduLcpot5C/uwcLp7C7kcJ7w4t/xwQdfBEcdyNcXTkoxi93Gae8PxN8TQJH7TcoeQC4QTARPhA/y
wZYfaFn59uz4+RjnS6/0lUqxHuifqLd5U/ckxwSZ97tHTSks4kTj+bfE9/US7M+/RbwN5GevJcRISh1Xa61nFZuP7PpYuwKzFQou4bIE71xUUtVwJAvA7/CBTu3vgh3+
AwUhxMWe4wzGS3Pn1zZYiZ7MiNTxByMwHKIWoM5K5wEUikbQLhTPvRwufGIPDf6J4qgIr5asJcJSXEunRJjhMDstfXN3guAoQ2zXtohnOXMLmy3o0b9YiLkgTbQULT/I
Eu9MNvW/E8Nj7EeF1wAUFuvFhQttzk9U76kNHuqGjoFt1712eKVRvurBx7MlXULEY5gcrXlnDl40jgdlQgwJT1IMxjGCOZcOUi5KCtgTEVsMa6oLzEE2KaUqro62jVhE
6fdNBVRJ4UPl69wnPbZVFmJbt5GyhXSuzchejGIzh2EW3CU5HUPgc7gu35DOJ//0H1FPZJQVF1D9zhDTUlr0wqn8vAAiZQIsqbzl9lVirNVH7URkJ1Ihij0axHYvf4jF
pR6tItVv/VGrO0aK+bpdbImx5h3/9vZS1QC+bqr0eGxYvGa5Aj9GZ/fnHTfD/gTQEs1+66C7NhE3mr7268pXw59z6HjnNpxnuO7qAp7ihXFoyCQpzucjAyqVtZiiNIT9
m63PXGohu9vAsNUGwewhjmVIhrVlydFPSMM7IWhg9SAZ5aUv6yeOzJ4KkpYQ9Rk1bDLlC+LRUO6a+8x2vi2hbmjIJCnO5yMDKpW1mKI0hP1GRJy/5VttYASdM01e9m9L
28ZSjB/UvlvkRwPrjI2/XEGFl4oFiWLDRrG85lD6w+JH8vIrlZKeLhvb9CI9ZrUnlQMMB88Bdbjrl5XtSpMosVc/AVxctrY1fjn18xig45vHWebdlND4kHqJ0mURTDEn
X9/LrsORNG7lFcJ7o1PBo/xDYjvEWJUyhai5mO51mlA7sgIYL0u3RSw8AgCjlkjGz+lt9UTCTRaO83oXdfkZ5cKOZ9t6l5dVjGKrqaqxdOLpq57bVFPn5gh8VmCi20tg
/U3DlLc+GWpkYOdJJe5tIpik6yI2yKT5JJu/I6pZy/4jfHQS7pOp90hhpyMXqI6MytV7J4Tnh4CO/JZGYmsYkpQs2bNh8CGRwj6wiEDW9q7EvRJ7zeoKQW0BCD+XxWsG
BcNy0xL5JpHhqyY1MhBRz8EzXqWTpoBE78SFPVHAZJ3qVMuvqww7/0wEPdYT2qaM51MH6XheNbUCh7iSfsbyKIQ5OAMZGu1PXwE3ZuhnvBMr+7wCHJcY4wnV83O22pcp
AjgtXFG+3/hMM6Sf5Hks13PoysZ3/qmqvOsFy3B45DUgqggeyQr/JAd1Y7tiS5JNOp6EJ5g+sI857RXM7XNThp0f1K5WGsoic33GTk6bEk6U/5xZqMdNKEeFh7GcjcNX
6cOGhmkiL+Xce2+K1LDBZAa0IiX5ZfbcbvqG/jNsJ/eTkhr28EoEUOAvwUZZgGTsITjdrBI471zN4n4QizBAOlPPMoE+JC+RKTmShngD89YMNBIjpXvnivun+LAmsUoR
cdDSKLuR4aVAOo9U0802UM5o0yoOX21rFoAz9lX6ZykMGNyym0LLHNyd0xXidjO+csC+eObxaNOznZGzlwaC78ps7dFXzx3g+BCSkqwDCv9syDVEqekfRfq2Esjq1RLw
/ENiO8RYlTKFqLmY7nWaUF9Ny68hK31YtVIq9oEtWiD2wH6FK0/zVgiwkenzF3Euyg1OgY3CczwmDCj58dt9JyY9TVX72NKoARETZ6c0g0r9Ua5ilyOEgo4ajGgxJpiE
11oVQGlldJkgWnZd86MRemVVwOzj1W17lwC+D2+W/dvTNj2t/Ir3RlbQC67ncZIlWeIs6Xn2kgrgNEKJlPw08DCKh14U9eNj2pb4IN5KWpA617A7rzX0zbTbYg/R/ue6
OhxGuzoO5EaAAGKM1xzfkhfegx3qDUOyw5bmyAms6Upz7EsrjV7VaHsw8Fz5VXkmBO8A7Q6r4k6Nt4XxRNiLYtve614njCOuSpTqM0VQxQNFwDDSjbkANjNkAagKllhm
kA5xFJCWWe4aMG4S2ZuE6xWvkFa3cp1qYbC9qXoQLKz94pAhQlrQMYsnPt7fuSfcBEBnJmy99AlZfuGJjjPGQjGeE4qypHDDPfomtLjKfsYBZWihmvYNCcxV4A1rQq9q
nZT4GXsp3UYAb6vB15Pm1uVEhH5lc9ua6X/Bm+t+osrg8es9GPj1GwPx3v4KyGqyNiZhAqCzVGR82tB6Z6nrCmGtgmoEovnzrF16OGBvkbyLdTyBfIKtswcVR9WzdMw6
kzXF8wmw8sA212QHXB+XZQMihk2UIadtYJy6iOd1O6mCo4daMIsDrB67DWyUOeJRa/o1griyBvZelU4wG0MuQh22H5Sqgo4OjrY+/+18qfGKEApLj/fHZ0l/yb+g/IOY
3qPeLlSZGvJ42BNmpjiLei+PivEhNNjUs9hMSGdymDidTnRlkanO42hahFTS/A1+s1xb5YFkAyc9ukTaXnchYeH6KnvxBC5kmgk6lF3xnxXDbMmLPlOAQGCKTufGtjR0
FAdBZm0CGneaaNAZUy7O71fya3Gk1oKvQJ6CZ7FR76DEz6YnvPZYA/Vn3oEz3Uk5z+AXC6nd3optgusPn7ZdAt+Xax1ojhEtbIOOIGunZ6wUB0FmbQIad5po0BlTLs7v
TYIyuLQcSn5n6epr9A2bPRDrIqT60fT8uE7Tp4TwYsbell3o7CZ67yld5A8Q0MvAAoUo+9/25DccoobSyRIdKbg/lqiiApd+W5VoFk2XnuIOzy29RjlZN07B32sCgMzB
D7sgTV2C57hgQm92rjMHhcMUyRZmOarpyKsEji7qynfWf95v1ibKBafoLTXeKX92ppkjpIi0KwOB7BcFvsER/dy9EgkKFov7ppSePnO6oKQ4H2Kp7K+pe5Ulhh2rQpjK
fVTLOMSERDnzHWfbyjtLolv4f9tQXU+H4W2zK2rR45151XPZyUyW97weMJrD4fLZwWYxk6BoIAxoDE2i2xAmk0NzAVENcbgJ1mZJUniNLCAHHcEupfcQAWx6Kfvbj9OX
QL/9/qq3z+xN3OVyonBcHfn4/rufPFJWQpN9Vqd8bLrLqub4uRNYdV92crKtqDnb92IBxL2uOaPSxWnd9WJRzsQqYwV0dNxz0PzYXnp4R8pgSJh98ouG5/usFQM7OMNu
Pp1dlAhfLievUGN+3amkckbVLvdhqkaqTcKPImA+5rw/IVG5GpV/w5y3h9anDpbsnNlBQs25VIMYOPIYLwxhzdjl0VJ12FsinnlWC3IjoLLmF3X0DNhFZKndm7KzUAvH
HmDeyngWlW4+KIRMKK0b5RolSvmhgpB1dKbGqZcjDCKgpKqA+mEWFXa7ndAv57e4rQWSTcJrhWP2RN4GEmqY/9UnNlLIzwdkSwoMY9YVvIqsjAu1ujl2Alab79G+QhAr
uPfMsuc3TGtChZqbFaIeLzDND9IUe5wgawvGByIZcsBMi4hZ157wLoi+hIPg0FxkQe0bbSa7PyBMKcKc/q/QeXxAX5JPWGEzrD/W+RU4uCRax0fclEy8jLi4mRN5vwp0
3ZUHM9RNAzXOnQRQPIJvcPFXH7VbbyL7X52TKNRzrmiVOaHDHo2CnOOdxEwODPTyFe8lOKOc4mJ4ll6aacRqrlYtAlSyXhDJ1OQhj1YKHpcGO1zOyYXgLQZe1WJ/MKeJ
K3WvgCskBQoxm5jAK6DVeDldOdzFOYxghvkCMgRTFxzpZvC/HRqVUxv0hUYJ/Pq3zq5zGJASFmizkXxRYyhIsF5FlyFPamuzFoSp+Sb6mlmtBZJNwmuFY/ZE3gYSapj/
Lud2nuE+g10FU5BMApoWK0YXa99/dYkBBUJXTruMt3LcXyoyreEVdZ12EdXnJ6IZdlHPgiHCyRHcqMwaTeFEyNnPdh2L+Gm7b0aVZMQM280hgu/a5VFoo4WOp7awN6q4
osuYW9XxUBH9XJt2Pzvk4AOnEEQdcnUYRJLzmhyvvDGAkWxR0btPDQWu6Irx9MH6TdboDcaP8nkREWZF4t2TgGVR9vPIsGCdYKHAOno4Zu91bgt8cyddkUgC4E+9S9P2
dTwHlN5MK7eudTyPvIRIzIr6GwF0iqSzVdwWMSBjCAOeBVsifyaMwGGheLfLvm2EubZ2O3niSF0IP3tnV7APHwt6w6CQv0P3IBRbPY+aXpHXyyWsqc58PriHFxmYmuHG
9fpfHDyYiJC8kBCkkin31u2eKvxL1oiNQCgkJWnyievzbVVieLn3yovL+DjOh8J61JdxkSPww2Y+djz/GdfmU4ALzI5pQ1cfKkXYUhiCmyH/T29m/oouokg/pLxLcFdb
zAT6vtWHz4wxCFHd7raKadNuXfmZVFTolofWA4KgbSibAa6RJwHx5kG4kzwqno72f94bQ2vWfPfaYtiPvxCp6dUc85FKIwRH/0EhJpqOOh2fJXwDfCW++gHLBv5pF10s
5DFgsd7UpFzSgGDJZPGylSyI+ZN/EGfdBA/1ms7aRbnHvFT0MebXcpkLvrivzLTquFKM+uwY/zCnfeGjrn4ePtdnFdPhAFTiIdDs7iSaw3U575HuCWo8sH9Z3cagdDAb
wfk9VU5Us+IBBZ27hJJhKzu0MZMlMhaYZdOYNnu7NA5+tH9kQt+yx8mtAw/zr42LWVFAy+Ij1w3a3Z/GAtXtn+cKaXkWHQBkKQGXPS8xDUoINplC9zlPwK59SNNdSLvu
ezUplJyzCDh+Me67f4axy2mIO7Tlan130xaRp3Q2FU2RQPzzzY4MiyM21KsHp1NtWJBHcAwa424uAmDvKbQqKSd0RvlkkWYDnKRTvpu4ZHyiIiuIlqT5DpyMhG83ImZB
NSNoODelQ4W6NzWqpGVgUekuKUvPl91h5INtKHQOfdxUQC3m6uPPzCmycrp8OzwJ2M1JYPoZmRRW0eRZq94u+lA/40riVnz2p/Giah1Eg4OUGMA/I+vREWt7fyuv8atA
uICYQWhiRF3dKhcLw5mJzOmu6na4Pkm1sLgdnxR8Bf6J+HYikOB/Amxu4OAEzX/3mD9iEwfnolhxE30HOW9PDulG97qmRx3YVxreUxfZXOZw6BFYBVW69cUgLDlAvVhW
uT9ybTFZVxBezO4ogumP5feI+Q0gCz6Knu/GT09Q/Fngl9ICWD3tlvYBsvYjngO6ngfifBq4mPZgszrtzxdF9oryXj/LZM8UmCcMURzgMywj8XapZ60wXcS/mH7356O8
OKlyalwBV1CrUcs/zFldandJufVkyEeAG3Ss7SZKVmOgWd7He/w1KrgMb/8zWm/wrEoeSIrRHmqA2C8hy40IrIhZ9wgoHZDpK8WzIEy1sqZEoYL5n53EGBFrg7waUa4p
S9UHj/wuDjwTzkYr0E8b4gEmVLodX2Qhahxp9CZsILyaOXpIngwqj2sMcj5dPdbIo/ZdRnsV/BbKG7shtNNcVph+dDyrn1i8AQmg/r2PaqcUlYfCI1iODoMTZvJCrCkh
QD2mxhE/53FPyKgc9imXxNWUdg7nBUYsmFggq7h5CilpmnRQv31uCnFBvRuUj/yS+H4br099SVNngJx8u13m86jrjw8uiVZ47mBdti2RhQApLD1/SYhYYezWhfxLfcYn
PoxadgOa27AT9/lZcSNmRzeVupLuXAciJA5mqL6mIyFXCRybDxRCNMhj2wtW9+9ZvarsjM7fPiUQboG3SBqUZMeBG0hUoHdmFHoYK/wG/wmulMOgAYhNhNo2IYVaoDYh
rEV4oWo7UtCrNgYwhhG/0+PHWesUHWa4V5nTXuI/a1TBbl/lgZZ5tuKoXbhcNCn7T+nor7TGNW7/0j0Cg2DBUcVBn1c3zuJUlktDH3JJZH7YsOfaObjrYlF66d5iwVYV
J9YA/rjilrVSdyXBEbSILvYth2+iDjUM/3n4Vwb3wU6gjo48xCJojbKCiOOTs1lxYiZsEWL4oy9m8M4GkagFiaTup7r85x/0AHOinMkSTBiFDJtoiO7MIsOJiES25/pE
ycspSyfQz1/ZwSALm467gbFY5qrWk9GrzbB9GQJUQUxkSSMTpVVjdwMC5HIfPyrRF6oQggjXbJSyItwrH6KLjJ6X+AuAEOV4wgWXxUDV7UQ8f8GXBSoggavfVfrJligG
/eM7A20bxq9cJkX5/Ws2RINYD+i7dSa/vY2Fuj+jOSoKTw9sVSD4XHWcseNEXeGsJoNfvpsRhzB7K0V8QGLVF3K6G+QmcR07hlZEI/P7HxmVxJzS/TjY/sWRKmFgqfwS
M86v6EtTY3ljPYLkCNz2PSMUfUAjxsgpwadL5xJ9/qogRj0ip1GCTUMZyzXgb2n6YmJ/GbxJwpmrgL6tKQy6fBAs3/d0mhHdO9KFY5P6NX6VwsPRQTZVudb4YrA26yAW
Nlw4TBrpZH/udnQlbiyHSYGGV5FFKjPsSTdus+XOqGldFJn9j/XuZWj3JGL5jIB5znggpIQJm+D5pV0Fv4JCboMeesrJjBo9OLJPyqm38ZAEPJLmUgawjNqX36cwuXEq
tUqfv1Np1Et6djMRcGANXwjLztOUOEDf/UutdC5I2aZY28g6vcKVCYeg+OlYHSrVnUlD+YegJdja/POQY1AOQ+Y+/9tbxUyI/NQvewiTUJw8KFki9jm1B6gGdhUJfpJp
orcryCloFigeY+4xVsu8Z5POWUK+ikvkoWaYSQI6faAqrIr38Gc37Uomu85x2YVwpal93RKzf1yT7ysMgO8Ap6FMcIEHfmV0pQ4Hj1tKiE6XwWcAF4Y/HrDYKJaZdAtq
paxE19BuajKk8dnVY17/a6zZjRn8x7VJFdI/n3SXT6Jtoyls94diL4HR9muTv8Lf9FBvZ2L5F9aISvOx20ssKD7jnoYoa0A2LHPYKRrfqCg/fICR1o73zoyWUDXw3VPw
ezUplJyzCDh+Me67f4axyyqA7KmHsyoQHrgjwoWuNMWo+/CT1ak3527bHBMaZRI9guMJbq99akOlUkm/sppZ52mbnu3kS/CsFHQR+AJ+5rc4dpmpf9LRHA/v1CgRRtL+
gbIggBs0lGeCTQCYe3GQOgUSDXKdrzumRJIY2FlfVnJCp0f0GcHScPX59YyEcCKpY1kc3VFmLnHkAVBLXhxN6AKeozaBrwhPFCBXdaP3konlZoP0oDL1yl6X02xeab4i
momYUPY4xfCTPyDwoTqFsI85SKvgSYRRB2gaQpkrPMf1aP2z06t5RIlZKrfdAcE9PFVGTfICdjHeyKM/zyugyIjxZk3gleU8OkTfg/DduyGOLpZUR8qm0RiPfzXCshjW
ZIXPgce8kFqAubiBWIvpX+ZBLROT+ceUOVmLqQtRoj931YcLbR5oa3wm6Q9s4sZClDbV9VKX0L2CQOKFi5H4y/vNtO0WDNjAYLkg23ZoFgYYYqOVEnPsvKhXIgyg8/rw
9rQBHXKIV1aS5ckOR08nNz8gAJpy22Xgk3ZFR5HTZisbX7Crr1onnh3j061iuTDndgWHs7HLmhxcB5x9V8XitXVj1RSFj5s4wBZzWj6z+R9cjL3fyizg+5K6cxpc+Uw8
MuEDEb97NJch3gbPCDnRWMi1L14zFd/BPmPwQn75DIatyQnOGqcnim0xXQV5DAfLdBFApDig7dlvf9JuhRnXFBcBnon7ZiP+C+Pn8cIbRbjsFQLHxn53gJNP/34qDtAQ
MbvwUppJ4RMcbZ1Rxc1skMi1L14zFd/BPmPwQn75DIatyQnOGqcnim0xXQV5DAfL2U4Lx1QcFg572690s2bBKOyXWGjsPLj4qZ4Xi8pYfDy2ybekvkMQ415iw5WL22w+
+jbikJTDv89eeZJoEz6kox1PO4x26VO66sW5RMBX5HTz3t3K6lJLPrvZaTxIZh5IpKm2jGp+DTZmkGydidDn5+esaTSPQ0nHaFaEbN3DNVyLATc1c98B7cTzThzla5xi
rPVJmz13lJrVtcaXDz5EGR8Z79//fUo8NPmm7OolpwPBvpHgtn/5fQ6ovggeHSile/7JZZA8F37vBUjB+UHNQeesaTSPQ0nHaFaEbN3DNVyLATc1c98B7cTzThzla5xi
O8mX8ekiiyOXaMBBgtCDMXVj1RSFj5s4wBZzWj6z+R+LRdJjwxWwkqIqIWen7d7SrzljGmeVe6EY4YD4XzxrraKZA/wOlCBWhCwNrDTT1lbCjHtMUWGtwA2hXdFBn6fC
20BRQdEcLdVt+RCvWUTim9dBvPl0tHQ2WOG5pZc46VgXivnxwVRtLcOw7KIPPEh8yLUvXjMV38E+Y/BCfvkMhjSIwJH9ZVmBSlX7/+HVOk7vO/OT0IjLfI4m1SVRPXQe
G1+wq69aJ54d49OtYrkw54iS+q2OOXhuOwJ1w2FwPMrIgm48gcLA9dSTDK03qkYWG1+wq69aJ54d49OtYrkw5/DSLglawiWIAmqtadhlhDxvTvUR/l3NAzH95S6Jeeu9
WKvjRIU7ap61NU810Q9B8LWDIyfuMIzvmbtQEkXqKW/04nS2XgF5r07M2qO7lEfxWKvjRIU7ap61NU810Q9B8EhBSzvMfiy03MKgjvXMmszhuz/5gMvT1cSc6CyNtPUF
XCoQCG8UZyuTbQRTNzvZy7FACX3z4oaApdVqcNsRIYRiDRvSMRUdOy3G4tIwtiQlUVfsPsYsEXRaIOFFRlKzTzOzwayX6AlsyMP9RSNg8HAHyGJsA5FiWJJP2CPchFPq
N/6dZfd04H3/P8sCCmyH9RoJo2OVdS/fbBRTTGTn0bzA7hZrcJGsgqWE4mHwsedkRReApJd2FqhijpH5FwSzevS87JinVeBNTs4XvHiFsJj9T4ghHWsSgdWv6Kt/m5Vd
xO9pzTPydFTwHa1H9Pm/oY/7WLoKM/iEkJpgCigshLbePXbrmhID2+9Rm1xJTmk4chrDlCBQeTn+cGc2WiNqc5t7j/NJFLNinTmXaz6TxCR67XyxTT2UeMy8vslQAfik
jKzLj0rDJSDKFEy5QFb3TQuVw3pzZBfDMr4+g8uePLtdeHsyTU5IFKQoBM33MA6jnzik1nusnalTVjHXrYX9OPSH8Vmo95bbN0HsShXdG86ZAKINNp3T3ZOhDtSyhxEW
Hxnv3/99Sjw0+abs6iWnA9YRHt77bf4CaLHyfz1NIhxiRiFn9l7UvGQl1F5vswpUYuGjbHMLjEp1uCl4p0I8TNCPIVveirme0TuadnQ6PW8m8vaf646NvvapjbyFdoAB
nT3w0cjKg/Wv5W/QDce76YA10+KHN8z4S1i3VAPexnvF5475B0wsm9yfT1UCafPiIfnmN+cVLqGDtwSMf9pyq9xzNBYM1Lzzgm021lhnjqIJDxVyEuSHFaI2UYhUgFFs
4dvGAIQkkwZuG/twr0wFRLE34RysrubRQFcwOjWMKOz1W4AYr5J4/hkM0gvfMtI1ZkkGzoHQvyFduVgn48tmDMw19TaT/g4P/BvG4cXj3lIBHgHGmJwFJxK9pqg3UhQC
VW0cjX5lbwqZpQb5zua6GZl5BGDTQN4LC8jgLRXOaME3vRCgOORQHfaYawqRQ1DPCJO2eHHKQRfQIGz4Ftl9r8NDPmyxAlzM2MtzUXGNyK7SMIdS0lwaQs+r7ON9ESqw
3OHwMErcaxa80GVyxXKy3O7AN8HzHMtlpz/Y/ZXPx6gQO3EUImvDNZBVAjJ5rC9+FwGeiftmI/4L4+fxwhtFuOTxj2mkraKD85a63foF4gHOC6kc/Wojlm14WOMPcALp
rYNugg0OZHRJ0OE4BZGlV3vqRhiFtFixM/THXVK3PabdP4TOG63IZJwgnnkphsZB0AkpPlvzv9T9iIl8PkAwNWhwqoNZYtGeMhcK5i151coB1nvlcnGk2KJd7JXO1p1U
bRxyUNq8UE+HW9PW+rS7AZKOD93Yv+D7B3R8vb5r7MUPvk2Az7MSOjHyMGOiOqPw+5w/q6ksg/yNR3GrQpafAez2MQMLRRkRzBsKcIN8XjmANdPihzfM+EtYt1QD3sZ7
PToFj7wHCL/1cwScfpVIa1NRUKA91JXej87w8UpsZbvY8QbdKsCF5+zXvYBV6zNU//CnG/71OApH6EmZn/m/QzENCFJGWccQ/MUKqeEhkrOUx6xy3K5jGbdwxlzmTMZ2
ePTysSp91AT6yfoHRTgBa4Vja9MAWp0VMLzPP0BZPQEfGe/f/31KPDT5puzqJacDY5e7dc9cUf8H7NoRDl+03kQzGw76DZhlQclV4wPtlkUxFy/FZY1l5riCSye78Y14
YdsoUF6PqU/+m/n04I3YzR5rsXET5uIEpiBJuzCxKy2OFrcVtiAJccq4tC2WxMvpkJIncPsH+T+ujSnVWugfJg2q/GWE6ABBuENbJwVKslgj8XapZ60wXcS/mH7356O8
OKlyalwBV1CrUcs/zFldandJufVkyEeAG3Ss7SZKVmO5SckJE44ze/uzWsL54+RVGS4cxUOY9rwhe6S6Q0j7pb+YadlACtffQKw7bNQPQJRUNHXPEZmiZo21v2oKmCOz
n+EIj4CDKvxl7RccgEUGs8wq+mKQZp8K5+JcJV4k7jcZ0V/HFTcMRiCoUo6XdkTa2JEH70w688/b8xsparkSpRXNxhaqfrXlvfh+zbvkbU6u/9ArBQWGB6YgUW04cd2v
xthiHOR0eNRhkMps5WcTG+iDurJ6ufAf0A0cxr6KeashMOux1zwTkm39wR9jEhXc4ssm7OJeQ8iYTi+oWiG06YQ8zvozZcIOYb+Ptm2ihmbiyybs4l5DyJhOL6haIbTp
5Fxwq0RWGQjwb7cLf4OcXqT/KdjP7TByw3oET198vD4wxb6YC7XUiyBDRtQ4FUPSIXHf/vjQVRiDeYGXBMr9lDdQ4e0KAlyKqVO6Aa5vPOqUr9L72QAhRMfjbBWXQ8MW
gpX9M++Fx5Aq4mHi8K6hQCGFPvzREzDYRdFXq1rp8orZd1wydoxoHLb0FG93q2ukyY/5+vr5uepEhywxQNnb20CfRKfmkZ6LsobI92SlG0JyVeoKep8/ak9z5VOsWc3/
L4P2vdp2AugNelRogsYxCa/M2r84wlw5bk4UGZSYuM7ZN6mNE5vryY9k7y5VvwpSgE4WCevMCVeYHyfw8VKPD4kIqhrdCUO63+5fFBBTCokxpjd65FGXTqrW3Au4e/2a
EuzmOM+htRk4dtQKCFopxtNQh43/wXeG+mlf25xexk6SOuWLdTjqojSTmiSVuTgzmX/1ToY4Se3bRIOW+v2XeI1pz/usQT3FlShz/ENcvpoed32BS7PggG4NgB7g/5RY
4dvGAIQkkwZuG/twr0wFROkpYdvUDWRfSEtuOkWh1S0kYBgy4TR0f7/Ziu9JcJRdFwGeiftmI/4L4+fxwhtFuA/+/Nh+rbYvanwIFneVgT/P0DoE+3o8V2V54dyJnMrx
iQsmZc+A+c+snOgzD+BzkVFX7D7GLBF0WiDhRUZSs08MHV2TrtVW7YgWLUsu1cJtSHMKhl+BH+OnqpejLJb9owf1CmnEIb6mZVJpTlakkId+o5UD/F1jZF/lVWLPaMd6
S94ok0ZRZA1E//NfExEA+CB/fuklHldwgCD/FbT0HTTIV+JfDRerT+X3WK6irfpf9KjFNeNuOynVeHTQ843k6Df0fgQN0MksKI5elrI4q4wfGe/f/31KPDT5puzqJacD
IOStNH4rCQprz225o3Esh3HaarrQfujXO7ryewuNEO0Pv7lBIkrsrvdlfYBd628cspw+vaujQGXWLezs77CAvyt+pHVj8q8nMSQHLa2Q4IgXs//o/YI5biSpjHZ7wihU
NUNjdA9m+YhufIykDBI7LSfWAP644pa1UnclwRG0iC7su5vR/JHfpHnWgbkpYuLHo4MXQYoE0+Vlg2fVykp47je5Z7TbXKvu767RoFMWtZdR+E3RpZPSOvl1vyiEPCpr
S94ok0ZRZA1E//NfExEA+LknI4JFavZ4wgyfbhOzvplcpbRd+rnPNwLvZnhmNe1wWgfMKrp4uZLXMelnEXOT0iayprqujGPQDRI/DQZa/N0PKb7gZyHDFliyPMFbcY7S
tvMkQTEmGi0z5papmqfC1E5Gw2LlEfUGn6gdvj9+Yyj1aBTfrnP+8UBgyY5bnovYFwGeiftmI/4L4+fxwhtFuJaHTBUwUlZF6bj05oIxpujkKP9+jXSRjNDmGAUjtAfk
ldgNEnTFbMgmFPudftN4y8dz4DqoL0P0ah3D/pPtaUAXAZ6J+2Yj/gvj5/HCG0W4/DXvyj4AiA9hyqDXHGX3q/HkUjb5yEWKcs9SzPGs2K7ItS9eMxXfwT5j8EJ++QyG
WEyWW4VB/+YmGXpWxpPuIHVAF3S4OJFuC2UwgGcazEv1O4PI74obAN/40hwyCHHX7QHZcngOBJKbnO+hOpldxVz2Vu/HNeMXOw0q7EjxCEssNWBtE4IlXnl+aUkfw/vR
CjYpTsANR5877614ImWdODMTRvQwEj5VS8w4XsRWZxNyRFhv5ZLGu+r4U8IHzxYrAJUWIn3LXAwnGb0b/ZcprSt/BCIpSV/2zRXZ8KMCBJ66pV/1wTfoYv58YDDoPRyO
pCfc3RJaV53HpkNA14BNWVIaaX3kMgR4tnNADuoRMZv/9QCkMuTcqV4MTqCuyGqaKceK4mwAxoofdoHzNhlqI6COjjzEImiNsoKI45OzWXFiJmwRYvijL2bwzgaRqAWJ
pO6nuvznH/QAc6KcyRJMGFd+UedusNbd+CQNNQE8xKsrymdMh25n3U30GTApN1MWMQ0IUkZZxxD8xQqp4SGSs5THrHLcrmMZt3DGXOZMxnZZa7Edw2Dids5LIOe8qPY5
hWNr0wBanRUwvM8/QFk9AR8Z79//fUo8NPmm7OolpwNjl7t1z1xR/wfs2hEOX7Te+XJQ0XAEjfy8kwwqYzcySdXKr/3xaO5Wy8Kuv63FhqaO7L6OiIS3jA/eMWrrtEbI
+91Z8vvSJLPKgRGtxr7EwpN+b4FS/ABQ9MaeqDG03DFWD5liNY0nAJ2jLxKzk6Kg4EFOFkOPKxbttB1K7caZ/g++TYDPsxI6MfIwY6I6o/A/IgOj0dQgjKit4S6fqDUI
ZbBtoSEzY4MBC2pPu8JcPlL6rQ3p/sPQuqJwPGbZZ76p0GoouX75kjsx/A8tvZE2I3W83crEShsbFvzkNdHFKmim5P2IlW8mG9LLnCZ9//SM9BcXviCvlGxUbYcdZUAA
SP4boCNzqSNhhcolHWtu3ONbMWwd7rB1H6M/E1ZrC2r0WZdIcRS2TVgX0vSMlVBSs+jJJnXy83rtPoUXRSGk8UWThPpy2h8QGQMia+GxbZ5ysDcD6YzqH1P+jf8Z0L7E
bUETruZKbFpDDf2roVy+bGqGdA620k6OhHIGypDJ8by1GONTDrHOFf4PYZGfsbGBYw/WrG+M0jiHUvKpmOsg6ci1L14zFd/BPmPwQn75DIZa92w4nmcV0K7t2qoxqBM+
SYukid1CuC5x8XSE2Ub3Jh8Z79//fUo8NPmm7OolpwONLhVW+GsmkRz0VAN1sWQ+t/Er43W52KLoX6FcF8+KRVlWbVZwZnTJVDfRe5kx0NpotVx1MLDzV4Co1CPUYmbH
JbmbAs8zlaMwNLipFetJlPnefNkDLu24v9nK4fpyZqeMzZU37PpFLajgqMr8EsDKsi9Fhl7fepBSa/FWt+5bnIaMKHEO5TNTS4kTb+Eq4d6kmUrsTmw1hXD9C4sUscam
Am8cyLjLTqhDOEgcd0e8bnfxqhbqrP7EMwSPicu5AiAJfIu/Yiusv0yfG1DMG4KfCO2CoMLelOubpihxFasT+pfGh4dhSdM5t4ubYwu6c12G+sZWXM+4FF7ShZcb2YDF
odwOoMLw7XRZdn8mx/78wJmQyKLAIKMHLCkzb7ploJIXAZ6J+2Yj/gvj5/HCG0W4954ZXrSGEBb+7kvP4D0G2lDPCRVRmFai7GV7E3WCFwEZe03JEJpBAOgZIYaXNL86
4ZAQm2hMmc5WEZ73sTqsNKPuevyUKKUdP5wVNYEygyIebkhjQfSE4H/ONyPHGL+OKHJQdwUQkj5WbOW+7Ba+DwzTBrV7cBy3g2PvKWdguHX1MK6fVE66QfU+Io2qKNsU
GppFIfmGui30K8Wbg/S0P+M3gBm9/rxBABzfizSxByvdB3uVWryzC8++VfBSGT701pGAXZRPbLgqIBFIyFnG/uOQCY+FoFvJMGMk+z31o7k/MAPqB47HhZaXfZ9oYWKE
ksfbida3aKF0B0dtb1pqPgvHT2qn2tarVm2ZPronYtpQo9/l3oSM/1Y1CLprIztcx+z6wrCtRNFhnPJIN+Yk0VNjTK65cn40qxTuLA8QLllHT2xNBk0HodxBIsltHYdZ
pLDXZ/iXXGCcLGXktG2LQiWIsVhg4TyHUKMh9RQOe7qsN1yoDKhpbACcsIXDDtN0ej6CtSZjjisBnm0lE7LP+SPd9/wIkWpkT/J65QxmrCAijyBBalafM9NLuiNhnmsm
OkRX6iW+aUgY9mO/HFrihWAHszZ7MVpMmjET5ucFNf/bI8AB5m2YBy8byFKA87EeW0fOXQMcJ2WNdEFFWfbr7QhLn4tBCftADTEz7c6sQd/ORf8rmpDfSvnwPRchRWwS
gkgWHHFLpm2iM1ULiZYDIlir40SFO2qetTVPNdEPQfDwcyU5T48Um8QnauPC6bE/v/CtzK4fOb+DdJwdO0DyjbpqMBSOKpyQUcgjLeugtF5kZbIIAucbPgGllk0BTWvR
FNM+E/RqIZu8EHh5jH/OPltHzl0DHCdljXRBRVn26+1tW7FyVCEuxTafz/bvpk1+/OzSIyyQpkw6zHlEdnUm5LJ0/QrDK5HaMdwnmy0pNkj+chh/dkYMGRkfTsOwNkFT
G1+wq69aJ54d49OtYrkw520yygLFeypZYIAy5S7xMJnItS9eMxXfwT5j8EJ++QyGqRzlYgEX1lYBSPBYkeEHYitKIBFXlRBGA6qVVjZtAcCh3A6gwvDtdFl2fybH/vzA
DOFLdy4sYRadF1bG4xPNlJS5wzUSTFdbHUIEbixPrjUYNrYfmxSsh9yY4sl5MEOJtNTLa6qf1QxwO1Q9/2IWglFX7D7GLBF0WiDhRUZSs0/CjDva+AwJk76QdwxdOWPd
SFbCDdPtV1TjOWgABrJB6mjrYGOrdFSMTrkIsM5zuZgfGe/f/31KPDT5puzqJacD/dX+vlwGt7G+Vte3n9Et52mh1/ZKlGeCSLsJaCO4Mee535sfg8cR0CuZ+51pa5Vz
UtbmmVUlbJ67P8LAaZCbuYZylOdxN4r7U7AvqtGhFbG13tRCUYtSiapLLPlk4hblEEpgAtiGRy0EScdb8cwacDjWQL6j96GNboRkpNavz/akWVGVDmRzFf0+zuK4H1RR
/5M2XQ5l45T9FA4d86aNpj2r6km7Q2bADtETGwpifQiRIHV1sR1AALENgNTIC25ntITvr8X8hQFk3x0CNm81qX/3TaNbT5FriW1a5F79XW6FzlbIQSQnFr3C7I66/Y27
7Yct2i4rQv0KVBSpkG/xMDODLYZM5DHkiMTevAPt6BJg5IJcVcbiqHTyZbAxqlnVVgVc7xRL54J4QIU/4mPXnLgBLJm+RWX2JvWpZnSaXLoBSTTwMu6Bt0hc0vVuhu4q
vRmaSIa0w4ktgDuKW2+dhyXmfgkIPxmGzBEPuxJGK3aSe2SjpoktYYnokSU+frE8PavqSbtDZsAO0RMbCmJ9CJEgdXWxHUAAsQ2A1MgLbme0hO+vxfyFAWTfHQI2bzWp
f/dNo1tPkWuJbVrkXv1dboXOVshBJCcWvcLsjrr9jbvuJGcfp8WWhPS3/upljCVkBspkmxYuajaWUWDrQtLcjIbhI9NEkSKuAbSUS9Bn9QQ7yWgwuV1haagx7KgXbQKE
v0JANQPQ6f8jB/OX4Y52fRggEYL91BBYBEPfKyMI2bd17T4OVcZvin03OnvckG9+GgmjY5V1L99sFFNMZOfRvNeTnvm1jq/EA2qflJW0q3iCEwrOzV9wKceXz2nyC3XW
22KCrcJv4/Bz/rtdk2WaO+BrUhlsaqH73JKg1oSGPR06KYPO6Drjub6Iu8gGHjben/5idKW60drnO/Shg5j8ZltqaLJXb73DRwdQSEKnTpZzFKeXdAMne0EwK7t6iwr/
BcC1XEksinneUTPeWY9M7EWdDOf2ngWgNVOPMn/ClHFImI10gUMAkfPyH/WBItAuziBrq+d6qi+bIHCKCc1ldHq4FD0EZJaw1RB+1v/T+No3kSoVFcejDehfx71AaY3W
b4pu76eYPbYevUfVVjGUAvkexpoAwHz6TZYOHk03WNko8dY1wNvJ2IqBfU+IIg81+R7GmgDAfPpNlg4eTTdY2Tr69bi8xyH/ATph7AP4WyDFyFBKh1c1WlQEHKZ4WWM1
JbDaR/vUSxjpBcJ6XeYWbIdR24KS0yPFGlavDKYRL8OGsxBUVdrCpiK7DUGRMFj+bbveRSnRu1owMGmsszz+2bFpZkqgN5+EG0IcMP6nGP8fGe/f/31KPDT5puzqJacD
iqn0eNN8sW7qrDH5ZEGOi4dR24KS0yPFGlavDKYRL8PspHLT6DeoRtfwckCKSWRMuBPdZjJLUuROae5tMZpLoAg2dDhpDiWeXVrvJzYIWqYmLsn8VH5l6QbPG38ywYVQ
fsTNGYzkUD/aD63lbb92zIA10+KHN8z4S1i3VAPexnvhUrOBQbaPn8ogI/hISesjn4OQ1QlEMiUS51ZFZVYgJI9jMzd7Ydndag3iP+4VOOzYMZN8WbIGCWZk7tiyDKhg
AbHmCkZ5sWY0sga/R+2KVLO3gUkWKE3NsPHO4uV9s9kWGUMf2Dx1ZHy7C8JPCKPouPJ3eLsa/upFRIShnjGbJFC71a/AYzOKa0NJPInKS/h/a4PdPTrrVcy7l4mrtrel
J94eY3uj7gOLtlba3/kVYCYuyfxUfmXpBs8bfzLBhVB+xM0ZjORQP9oPreVtv3bMgDXT4oc3zPhLWLdUA97Ge+FSs4FBto+fyiAj+EhJ6yOfg5DVCUQyJRLnVkVlViAk
kbbTjETnpduG4n+9WjmigLLuoJ5GW3GTR4h7MV5owNgZ3aB1LWsjR3KtL2bIZxu2TY3iXQdX1LvAGQLzbjqX7pAvwLyEOHhPSKqnDz1yyTxB6GJ8cg+XrM2xswNkhXCF
CJ3wWGnMTPkb4UmFSNSuGWsAeihc+xF4PFBeqorqf+CgU43791d5VsH6vF3+1RoauxcPpdWFkuJ+aAsAPIToGJl4THlHhGLLf8kaljuMFHaiJz4MMpGKeIhiepjRz4mq
MF2AodKUBi0d4kiJCbUizHx9RJLY9BZ4/90WfAJ7gbySuO+lBTxkt8ZKWGkeUjNpyJU8s6DH/JkUzQYL8Gj56qjrArWRrtwGZGTuOJQksZ2lQ7GMgY6KVSxeJ4z5CpDa
5ajw90Zatz627so2M3+DDip36BcxeSuC728wexmUPgA7lmQeNJg9br9Bnn6PMEDBb4pu76eYPbYevUfVVjGUAjxqj5TeJ8XjjfqeIzd0i/3hmlvNWiSMMMtjnyNM5h7F
KnfoFzF5K4LvbzB7GZQ+AH7Q0bdyNbZYs1YD/UaFKCsfGe/f/31KPDT5puzqJacDe3QGY0YSrR0avNa6rMsorLBZz2Rqvmy6Mb2JoSBhy8kd8JImk+sHQPKpYvFGEGeR
t/e9EmN7Cs2LYikC6+1zVQvOk1SGcklO4YoXWbztm1wfGe/f/31KPDT5puzqJacDMsV0CH4hU3vCOhdydvpgVeIJdGA9dyaiHh/bmYEhWhISh7BnbtMlo6LpBAytSA2v
W5VY02UDgFyLGX/OhUeMb43pWS+JjNdsC6ov7I/QRQjSDUwVSve7MQ3e610j/0aPHtv+TecTTw6/bsLFYXxrrOnnEjZGr2sb9l7Z3KJiLhEXaBbO7CwNIvyy+O5KT/jV
ZSkn/km/q4ClThKQpYIJBuKi2LceTNiBptSm3MJ0npDPyh2KXP/izOFMaSiEZMS+pLF0nKwVBiU6YlddW52BQw11a4grCfIbjjaz5tF0qusmj/XVeDvAHrsLsb/TgqSw
uYsKcnay+766lrxL6of6YoeYHcc+zw0skWvUjiqLBybjxccL1JsczA7tCxcRN7+oM2cGrDeTJe7hpTqBcog2RRWIB1G5IzwsYZG5SIo1Hiitdfd7J5o54T7ZAt2WnYiC
B76VDKQKy47OYeCI4FM8oG4D5FRm0JJJM5rZIxMrPJ4fQxs6jPMrd/aKOTYFDrqmbD21NhCYJHkHbmdwXPOhXbiI9nyNtXbyBRmApWa57HKTW0mYtZWlj0uvadfECXv5
1PkDfLcMO7iXHNaSpJHsRcUTerB+o5/g8NfJeRISEn7dVWckL8Nu3pVplAHg3uxGfnJ6eXtyoQVmncRXICBDCo2I5Z8gbbxVd0unZjVRg2H5K03dowVxwyJ5PVeM77MN
uR0CjQgqWKpXQUtvDDnCuwitwU/Xk5jdgG7HS4UHOWeKc5EFNLqpuNt8xx7V5d3eTD9k1z1eZ5bBLekLPQnCOUJQNxJ5qqJGIvmfIQWvNUWCKmEk5iCcRooyGOcUBWeZ
v+gGToFaEtif1w3wAQGkgtNcKgAMILRYaTGV4cKbHRm6or3RYGxtbQjKOisRvvFN52lepOGBgPa6DrxHHmrd5Q6RlC0NcZJuFXMODKlFbHj6M0li4v/vMAr1zvxZs8fc
EAKrTcPSQXpowDxSYK13aSW6VwHPd6LEe6i30vJzxjhP5bwy6ISUh0ZhPlODImMAkyv4F3vReBfOkeqSDaIsviJB/9Go9AeSBfl/5vFig/00f0jAGPcMVtW4lZxgsJBc
Dn1T7jgTkUzzBgwDf2RWOuFOkMyOzpdaLTWr7/n1kqDNMj3thXrXX+XsjSdm3mNW+i2wZboYYdMgAhCoWvkKWj1PV980eb4I5Oq7OFEikXs9iDZkZquzkFE227MiDWFH
Lru9lkdGWPtxRKlAhbNElsU30X34xUS/YkNQ6mPheji4ZYDtHJlRoW6D3dmtFxXfuqK90WBsbW0IyjorEb7xTedpXqThgYD2ug68Rx5q3eUOkZQtDXGSbhVzDgypRWx4
+jNJYuL/7zAK9c78WbPH3CS0kWQwEOQ9s++fqS/HJYba2habvGnSmf1Sai05xOhzpxRvIiw/ScgIUTZEdDNdFV3GtUhUu2zzCH/1r9l5b+aQggKWTglmuYaNYgx/I/GA
HsVftL3kjKQ6jCaIqzGe5AhEBAQxH6am+xUN7583e0PDj972QxizDcayFRUkWVhvvuY81iUey5dDwa96CP3XuzAtXE7u29Mx/AxGN4V/oDX1O2lYa+xnxSXFtovyHuDZ
QvOFHQ9xMt9WJNCUW+HB3rJQa8yORXbRPOzM7470nGqpMdoAbwZ1DGzdKMDbCXpUiWEZQK5LulQyhzNP2q4QkJmJeyTS6+5+mwSVvd5FvFKJGDxHbP6eLoLo2RMSlXtc
2IrAPasUl3yVzw1pALVvecluabrIfdrT2Ok8CiED+TLKj/GpWTI/qkx+24RL7uj2IPYrExlJYL8EN3PScCUov1XUrLZLe4yQFk4yl508P112vdCkpxTOUM9lYoZEfXhh
jyH3x2zw6FZWtlT9AoaDa+pw/rRylZ2639ZpoZKCYCLsuvxj8U3477Qgy5J3xoKrbKzP0Ri85GwrMvSNqBozBohUPNFNvn5YtVvolooI3nFXYWis+6idSIpqLx4vXoV4
dozaQ6lQgorQOIifg1A2rVzxsa3uozahgj61FwE2Sp/aD1fTeKzIDPO935hB4Z2lcz3OzeOTGZclMJBHDl+ti13cd+9tCAkOIh7HJEaZ64xPp75mlFZLDNBxxkX4pmJ5
f9Y/aX7c0dq+UIRr449xXPHyQTYJSG1TYTOkxhmQwckBCZ0Majlb/jmNSfVmP0JaCzaHSWsFr/rTwEYb3ciP5MsD50lIAhUY5j1Yp7YHQ0cOAVtcm2Nv4AVCkLSJQgCz
RgAkT8GzMh0Fn83U9h1a9KkwCjLVdup94mE4yW8yprqitBOpJViMYMkZSEN6r6tZzld8sjM9TzbPJP43FPcuDL1pjVNYE+6hPvoakSoyNX8QzAMvcYqKE6xKKyZn9Kya
8DbQIKGF1pc7av+NACxk8cgUvQi1fBP5Su/WmH2PUI1mhQtb8t+mYvM5a+hIxwEeFg9Cw6hbL3AzIspo32zmVvTn3XF40Kq3xjzW+2+JvAr0GUdce9JFsUIa/0kbegO8
KwT0XQZzUlFW0Ph3gi75NS1QPu7/cbuiOLEau3iv9fnmb0bLQvUTIZpHVcXznuPuJOgI1qtYPlFd5RyrvGKXKQJCfe6vjr3/hCz0CLnOarJv+or7A52weBIUvPBaon5l
n3+3KUcM4Eb0VkBdhMixbaAqrsffk3nFI3b1EN3Y5IgnzQkSSHtphpzQnD+jI3RRLmcGVQIKtOBOqZUQ8zffQgGP3CqGhexzxhHtCuk2VZHqIQvwFxawLkYzFOPBeGmk
szkygjwy4Otx8+973PL3tPnWXMpyp46Cgl/n39ivVPs2ITrIICyxT08sfDrItI3i6NWsi82ZbHeAM2Bj3Oeq7+2skF+C+a9CXFA03r/bohKaitwV10BUcBCh6VZOTrKp
giR1WAppcKd6NAActf1/eO5Jhqea4UTKOlW9fDr4bsEeGr4TnggugZ+4XcbPw5hnWsoTEDTXhkI8yulgVp992wUPov1zDRmvolNCYYFaZh1xfZpOtD4K7jzIZE6dQdV/
xZ4uUtKgUgWt2gJcs9xeJMnd0dV1VmVhvx6BPEKepJ13FSkIYl4Dtnx2pqwV8lRQ2rw37QnWrPcdXTUpH6gShxJgDWK2Hc4yblGRBiGvYZoQlzfYQYoS7uDXYg4ozfNt
cB5OYap+OkEqR7Yy50CfpnDXOjWjv10VK+0IV7zEu0BAUE+l5wVbRwQ87ivamnxt6IehNOE+LGwrnvnW4ns5ISOqC10NSIppitZvhKvIhPZ49i+KNO8zCQhctO9au25E
YYcOJUXljuEPed4c8Aktd0HYtISIes5uXZPkFDg5OAFn7UtkHg/FAzSjaNFY1g5rO7DhlueybJKk+vp6lfwCM/lYTBU59KFirisrG8KTQIQ6B8o48M8GDJzT5DGM7uq6
CQycyJ2hhMbsiOWGmK2V1pTrUdUeKq8W0hehSDbfEIUbNeoFapVG3JwNYz8rITi5joFbQ50zxYsP6euJwta2Wruc8RxPoCPDR6Rerc5tsbxmGFaCAWMdIPZ1rp0nZgsP
RX19gniO5FIwaSf2ljTvfT89S5o6Hiu2SriFNEzHkp9ePToGW6MN0HkI+4rhtPo5oRJzFF2jkMWwAr+YLgY2KRG8kWqJWcTH2Oy6GmBCv4NP1mE4rUaTqryqVFdAQiMA
Pws/HoWCzjoz2oSFI9+SThQpP/dQSd2nn2UKOCjotUmAB2+NGAM1778en2q0IMPSX7sEsop35zmGto/RamIp8jlFwaJI5JOQNbQCwah0gM+RxwPU0QQX2FwHrRaUoPa2
yJU8s6DH/JkUzQYL8Gj56hCD87D4xAZKO+7V6iptijwDCiCGpT7vCGg5w82Oit8FH77xJVugR1GlLpOV9ejwR04HUbQK6jmV/+LvuXsc846pV13utm1b+WqwYBouEsVm
calLfJq9mytfz00g4+hA9jxMPTuF1BtHZ8CU9S3T6S14iCFnAAQTiwMQ8utU5oi+8togy5bCoQLeFQmJZJNGociVPLOgx/yZFM0GC/Bo+eqNYN8fxL4JaVQBjDf30Wfy
vCsMnUK+Wt7MnahIwYUBA+TRGJBuxo+Kep4NOQ5JlqqL0XULqwiWvpC3VpM9RxaPG/+9MgOdNti/qdFZHsHNfiW6VwHPd6LEe6i30vJzxjgBZLyl7xBb3AVpd8PCWf0P
x1+jEAApJAKvSpIjEEQSpws0tYCdduVmltdx9FRcTN2juunyu5bbJjG01luRVo1vJbpXAc93osR7qLfS8nPGOI8WQpq8UT8tGX2M0mvAb+777+6Q2EAVrcum413tKwCp
zsgSN4GC0sr+wmaKvgvVtRySNiwKbcBCTQ+cWuPIQbxpa6Fl95Si042Z/t129MAF84WAWiHCYJ8bdsZR/cqhqnIzhyDtTJH+5SY00xFzhUpp2WpwOWEsGFFT/22TEoPF
6ErAQNUyspcQj5D1GajF9MiGaV6EvKuLVGQb+Og1/nufQUbiJYCyBbKmJaIjn8fwPt/PBVWtfK9PucpAEqtaV6CP54wpLZtRXJHuVzKY4vWhoiFXS2/S46Kt6nUNmDa4
zzoNf7F5ohpy6VNcUwrEMnU98A9Ir53febPC20KxmWzJBj/dEn+zL37mf9+fuUbzqhaUASgRSNm3XM5UuM9KJWh4wYDEJEmC9f6soEXtZFvjML4eW/eZ3GJShapjtWuA
5Jh2Vtt02g5StPoZmxYyUBS71m/8Bu/01WseMYks42DlSgO8eVV5wQSRLuADAXx+gQfMWdWqMYX9ctscpvC0UlUu7WNm4Qtt3rvGINJx4X46+7ukFpKL3BVisLsU2oXO
/t7gg4nusF4Som7xDNVI4FPIv9LMa5TfmhIRNAf/jvrAT0w70STYSu9FRRHNMOuXaZepReiES7CTMPjVWDf53fGJ1GR64bncUKT6tVy3PhuEgeZEzHH9bC5Aik+jtAvE
/KgjI5WnatXN2miykNGGwsArH0KXAXkQYrEidjJvUxPxyZT+8V53/j6U+2v6H8MxRPqCWvi+EjrbxGPd+Q45J69aEjbomeKAEONBdyYGwSYGHSeyiRNS68ISK1gIGybE
P0zzLluMLgJYBuk8DSrMAMxxjeUxWhcku+lT5DFRMMp98/1UJlwrRUGZ/XfvMZBbTFPHI2DMApof9gbgxFxO7vNQzSMLTGow6GRmn5uigj/giVA1+r0O02r3AhQDm8zp
vGj8frV+0nRPrMF8cOjXoe1r5cUeUhk4ypV80kv3/w9eYendhRYNQXP1gVsudbqP/jaSHtlfOUdLSzvp85O9mq+eXCnZDqUYxLNDHBHCGPN876G6FZMzWYUSIm30MhWS
rYaHFOyzcaR+98Pr6hodsvI40Px14WU4bBwHwneaJGR/fvAwi+dlQfwj30yI04LjZhNj1KVuIZQrDkrh4jYfFu8ZXeuTSBlwSwT0Zd5H6cdCZfUyO+Vbrj9MjfyFuI9d
Cra3rlLbtfd1FCmWimn5paaLAHzNAs+B17o+BeTE6XjcKi4f6+RVcAtQjBVjncMPa5cddgNzzmlgeiKOphq3gCCyNtS70t7KsA+9KU59RmkTX2o3q5noJkKlODZ6YXZA
uHzCrkNKx07oXr7XignY0GxuW0N+DnVrw7hGYpezyji9ixwlHjFMpdEUlwAzmS4J0la7sxkPQ8Py8CRi9WqKzuF4zLfYZ+ESuJ7+EnsKfleklgpnsvXJpAWHQT9VGP/z
r+upUehjDvg1dM2RHYommg6rT0Gi0FhHSrYWZ215CN1VA4Erw2IbBanXKOk/1+PIfOcctaXFDlFQcGEdfEAwEwaWeIsdeEP6hrcB9lB7W9BLDvPlmKbE5ic2M/ktNfw3
OtmkfJwG/2EuCSaRevPhpWcqLYLNbNeK5xhb9Paejs5AoGESxDCeA5pmVmd56fsoqVTSieJ17hRE8YMfge9baJ9thLUZVtLN24e4oorGTD4uVxgzXidzlG0qJbTtb471
UpF+crXDKtK2IQvyWMn/jbN3Uc++dw13UFOS6rQv+iJd9tURKknf5cUeCvo80ZcTr+1J818Ip4Qf/iI30tti8l1YVaiYjkI0hhLn6MVn/ZkWfkt93dFr4MEN035yS/86
iPNB/n6lVxu5SMEZxg5Xqgxqqb6zYOxeOCX+GJUFemYk/YXEnI6JwgSnLE2Fr3M8YE48bKA+OcBu+mGQ4R/GyPxgtJ+hb9jztJZSGaSErP0GG4RZV2Wvij4nJn+XIgHk
SbylZ0L7ffV2xgS8O8rJ69VfelNKiXeNkl0IP6JWfRBZWJt3CSo9hQi4b0EqvH5X4Q5vlf0DREIsDwvTk+KaYPM+vkcsDErE0evH13nrXjMs+eQpzcLdCW/7akqE2Ja4
Ck6lBgnL6gODI7PrXuDYcNWSM3hjZD0Nn5IpCvij13I6Qxe+nzKTdnf50CFA/izGEkZllzD1kPhzg9AVxeW/3U3mDYXbkzsmY2wWL149gjyjW3X/RwHgeM1hDoKE1bgr
vz57TC90N1FkkdqAa7YhZkA8vlTqlAJqGaT9+rbYaHRzQFbK8UjU2dLA++S8CKQLLWjz2kSiozuybniVKujRB3+PN7/M2cbshJzp6IyCXGH/G4IIaXMFp3rI2Fw1voo6
rVU9B4azaqv4TJNAcKxC98+M4i6JgBf82ir76efuu+Jh8pAdqDX/fGJoCgLrqwVxa2f71gAjd9IvfxgMK+jWbfEJLL36t70lEifW0viSXClDlncfc4/90MWZ0O9W5smz
J5PGk00UEYuVkNAva1upp3q0kxHHr2sfAbpZDGRjSOnVaYwnYN0CqwX+Ks2CCxG+8qNagmLeEWo6RuO6SEWLysL7WhenBtvh9E20kwknumdqEntYnUrh8MeaUZvmkj+0
CHcnHmbfWRCANczkAJSLlIqz/VSiWwhJjcEGgfHa6Yd0HdrstN63rWxLlMb52oqumX7nAugfAguChZPksi19+D3N385lokfY1YU82899Bff6jhnFXfZZ8Jnm2nFpKvxR
d3pJ8amfFCs1pMqU7/M5gnfdpBCxHyiGmM4oTA6tWgsc235cQoSTWoaZIxVxGGq9L4QCtPct0WVTjK7Hj30L7KgLn6MPdVOQo/WMhiQIElaRlbSgoNa03rnVF2EaUPBc
AgIQc62DXYPIw1mT+1a182Wrqp0tGUgqkTgJsvrGeTton9+KvtdMvtb8siFCRXHXI/BQ6C1yOAafNn0f+XkpneMPbktmePjw3nSiz2cS70IUb5JAWIlmvpI6FZnBXqYC
OibQ5fLKbSK/eJTn0/gSuNZ6Enys4vzh5m71uUGLM6nxlyCEgqx4/dVOhWNOCisb9b8gvZDMBAasph9OiY9HVMHYpdKMJNlKNXglKxjkvsEkcra1TwRWMhPXBmt2/Ybn
VfBrmPsF7zsAMAl+GcjpjRzzfdMIZpLUj0lefFeNbLzzqMFV8s3Q+4K7P++qKyvpQNwxX/4qF5mkRDaKvRtdYZFDnQ3ehMu43tP1G/dKBA1bxA3oLt9gHIexl/oLampV
EYIG0Uq3FAXekFF/l084K6XQOCMF55KAZMpNs8zHZ9C+vzQgvKPW7lPGfu/IQQAys1jklH4kkbu0sSNOc79JXLe4DymbSF8FjFqC/lBZRVlmR+YQjzHADBiEpNjgPbM+
7CBqv9udX0R+5hVyBjSR9zjJ5qWIGGI7La1J7qVMt4C1HrjaoapJGvfY0LzyBm10C6Yogp5fa/449/hH4ImISXSLv9yCB5fm4fTYiWcJSXjMCeGqbgbr98OZtno99VeS
2iYDdRv5xdnf1wMQchwUsvAzWsnBhDDuwdqzbeymPi4802M4j18ypDwPBZLnE2TSFgSb3qYFNKMOmNskJbJ9EktA8HB18nyxK66Hx9qDYSH0THXni81jVGbuv/2j4HPy
PcZ0ELqYDdaE4O0Gl4NcWbAsA2BaVcqzFXy4sABzztFF2SDOzLLhRA7qM5DIpKzI4/i+3qD5gwjKdXpB1U6jCkry9tA/X/jweWduYg7cIhseE/jIUiAeBVavw10LoaMR
WIpeLU++LOXKyhFsjretEvZqqZ+WD3tBUXuxionKle91nZJfLGs0BCWROHj56JqUFR3K/tbMyKmYWA/8HOzTOei2Z6grkvI1qUAXQ+E2oYHCGHh2h9Rlo3Y6pWRVBgc8
PERoLRIXuJJuX8bGWzKhgULYcG0cwFQKMJQIFA3agpAwWUIW3ModgDkwwSy9ntOM9jVddUBKKTE08rLvA6THgwXHl7BG7vshPzRCkisMARF/o+kX28Auydndm6jOZR45
LrmZboIZNKs/j8s/DyXClxyifUyHaa9YbgQa3H8c8TiEKZNfnJPoC0GczEyeV0zoQ0P4ZB6hZL1aXY4WXozXwYgGcLVzn84AusfWcwNgRZWLXhMrIyS22r3N1QuVoabT
+us7uZXnEXadhG2VuI9pzF2l6GJADnePq6wTFdkmszaIqF3soIrojq4tFe4RWVOD+NMR/DUI15lqXUeCtMG5DRceQX11iDDNY74oyPdbYQKsMFCBsCeL4wvzUX3lP53T
hFVMazZi5fcFeoBiogBcmgYKejlXtFY0AhbOejPd7/uvwXTJKm9g+XAJy5vQd1zxM3TL78YmRbQgCju76B0ggZ6CTy7QKhK+FtoWnduvBCgfpyeaVBdik0dNbGdHv1zl
sLLuWnVSN3yFzvjEI7PcHRGpaw7kFrs21kFxuNMbmzUOouJeT3/zdf1KkUDe6TcRt9HG+S2e5GcKeAatT2LojhozYdMx2tDAN+ia58gHDDY90OZmG087gCMQGzp9MHMu
/C9aw+oo+IGPAIZuWHAnsa/4mlUaIEqKUyxtHs2YS7qWaTniZyV/+OEGCKYrLBONPm1MT9RqKqBVrQ7rcksdgYrLj5bfn7+GC4T+HlCyNHigI5MYG4BQf8963Whq2Q8F
o/ERGpIA6JSGYG/qtOXQO8POX8x46P0xTfy3IKT3Kw2JazzFe6N2O13ZENwBuIIy9u9dv9fFYFcq/Asa8GEKu8kntbE4rTyv1YbFcmb5XG3gzimaT/+img8DgcGcb0ke
MjoXSCv3Ht122NvrVDxAtdEhS0DeckaY5bULpKLOPbSUGqSPg91rFwe9bi0y23pBeKti24DMctHNnjKuTUUQVrr8PufUHWBa2JPwE59EAQaUvUEGLvv0EqgTyPoZNvQS
kV8qLZIXxZrcmKysuQE/8e/sxdFnkN2VTYQcbQ3Rpd4mjhNUaIGkhYXV1iCQB/m58ch76jwkhOlBDQLmISwhQ7r8PufUHWBa2JPwE59EAQZ1ihB+AeszTFRcUCXlYt11
gHminanlGuHSwe6ovo4seKSznGVJtIad/4YNfcz8cgDv7MXRZ5DdlU2EHG0N0aXe80COwcg3hmdDOTKV8ZfK4xzbcbeofUFolt+KFjmqn6S6/D7n1B1gWtiT8BOfRAEG
dYoQfgHrM0xUXFAl5WLdda7/MPTuV+wjlu+V+qhwFZKZqN0A8nYkw8WO5BPiLwi5pJ7XGI4rLaDZCZSuXZQmGFLnZYx74aVHuDnOYri6Y426/D7n1B1gWtiT8BOfRAEG
ugDon8z9YPJXwP5t03fwNb+2J2DYV9VJFWHhJuOMHv/lsSQXXO/ipJNXeBoX2GeXcJsy7K8I38YTP9E//DHu2Lr8PufUHWBa2JPwE59EAQa+8XUXMI+vfYejwVWyo8Vs
eEWb1y3ROTAr/8Spy4SqjGdX+oqkrkdgMccR2vyY6BfG2bdBWKVPIw8hpeaEsccP7b0JguN10/zc3EAaVsqZW7LGqrzA0a3TXVNFwZ0SKAJiJ2BIM96nJ9zqHYcyuSMI
7vtCJPOuuhKGYTUMUrgboSgBZ59p93FG4fBVVtx0GA2M0jG95bUbwMCzVUJHZo1N6QGr0SMHa2RJcOvwF5oHYb2k3ikue0gaPSrchJsaLWY0V46anuPZBkOuz23p/+bv
ovLeMb4Je8gtEI4IUegMaF8zmMR76CXcIV94TLY+kySaS1005EtXrBoqXQqFdAsiDHDcTX8XoDadHI+yyf8Z5MoyShg3H/OgspaA42pwwllxnXlmcFaqIHTIemo5K5gP
YSMzPQdjfdEHakipTanpdJGnrmkA84TkSnQTPA3WD/otH73wj1QlW1qiS0E77BGHE5SFi450Nnc6go3cFYNm+rVB8U/HS5p+CujikcjzXYKnuIT/QU450nmNBTQhOYG3
r9FMTj4BlpqrvJyMLfWPf5gA5sjfx9Eflm6EfVjHMLyyadsFrhWaNuMVrKbTofAtbAAkfde32YoqI90dFQxVHn2aCtRqsW9xfe2WwZZdJ+OFYwW+foD/WvFT3eOtboX9
gOgyJdXQPceIbEclqi/PqO/B4HDywjmIa4RSELZ+BXu5NHVIBcry5zFge6TZNYSio54ehUJSrWeVFzcQ/VD0fe5OLTJzaB3vONC+Vf1SbMeA6DIl1dA9x4hsRyWqL8+o
V+goXDQEwbNWaJiUqja2n4DoMiXV0D3HiGxHJaovz6hMCi58vQcx4yUPHKIp1M2eiOJSfsAIXv6b4FiMxU/++SKFAb0TNEFHCRM/SPBH/02A6DIl1dA9x4hsRyWqL8+o
RMV8Wbms8qCsgtQImqOTKoDoMiXV0D3HiGxHJaovz6icRiemq2CvimPG3S91iQZBgOgyJdXQPceIbEclqi/PqN++iBpnEqDNhVKU2z+dreIcz0spPg9Xx8oZU3WtlpjM
CX/nF0Nj1RFkSXlmjb4QpTiLJOtKWwTHVxsTI5HdKoZtx+w69e1obHgbR+A1TJTCJZd2m5+U0HhqJ7J20BS01nCG/yhGnbhj/nMcyqHPqzGXmjkFwZLwugQzn1MCVqF1
Rw1e/OtUXRzfSfMn+rLCFlRHkcDwYl7mc52XBzANc/WBIgVmxK1m6pW5kN9/wGg+eRlp22F7QgOYPIKOjk+FDNHWWZ4i1pCSxS1mz96qk/HhFs1lzmXbiPfbLqC+h3MK
kU2Pwzh0bEo87UIuSkXK2eSAbk0Ukx++cAz3vMV/HpOPXJA8aHD8kcE4sDTJyX4bDvl3svaOsTUrmF7hzcDmdHmIcpAkFhFrOwUcCyWYeiwa1a18+O7gy6gxbsyH0pI9
XrrCDZIcHGLYDEl3UKCDXuf/Exwfs9vXEAFQLrLmMGXrxeAHOJK382vbs70aStr0ylKy+G5Y+kXrstr3BRfkV+o/VjD476MGn+f9qRJAcGLtR+GGtzKLV1i1uEwnMjoS
ScW+Bl9U6v1l4w1M421nXlI2L4NEOh22cqXi6uuk/BeV2qh3gPZ0xTotZscBJVZB1ynEI+XF3SnlUutX1lnLl3n54W4LJv6P4WmJoeAptnwo/vOvYMq97c0rMRLHMdP4
mMIozqg/ByZSsMh2jxmNLOIsl9qlXIwkM8y4nei5vml1QW7mFZwJeg5AsVzy/NK8eqrehIynDw3Po1eqoncPnQCpgt5FHru5iEdMKWKFd7j/ECjkjMbGzTdKb/rXusGv
BUoPIDmM1bFXndBwi68THS5dBrHw5U/SkRutL/IcP7cogX6Gn0+YqlC7Av0OdahsdJLUEdGm7kOlmdee2yK9HyS1kCVLguit0vQ1wMK44pmKzNt2QfVeAQVEqJv49/Wt
7/G9zWqRRRtavS/X8racHqablpSWzbW2S778l4f8U1gUT9dpXwPnuNn/Fb3E7IGnWANR7up35BPaj3IZ4wcvkYIkdVgKaXCnejQAHLX9f3g/gez755KbcRWfG/kYtfuO
1sAk+o8v5XtBmfY3SMAIfNixy45o8IpAoWrTG2aHQ6lj82ys6Yyrn0yjQFhOFWAq79CCkfkW9UBTSv7vYSj7RaqiKfatInjN4f8dRCxsWHJBb0TA7341Hzntzh4MtQAi
OYkTUoc9ZQ7NH5MvaN006voigaRxTfKr8esZx40zWLTtIArpvKivgZkiW5qUt5ZGThc4qqvRXloEq0it8t0eLm3wb9OJsbttDsBN5AROgP7KQpz96wlIQgvTbbQJqYe4
KS3ylyjBp1DPs69vmrzcVKMHr4KKxqKY4qrPhvP+FOodtGuzgquH7jF8JtqJFnioBAwY6RZN6jmdX1MTUxmPPWmyDT2ZGBXs44O/fZsUVSHLOHCk3YOvn6HB6K1PFxKU
l5o5BcGS8LoEM59TAlahdUcNXvzrVF0c30nzJ/qywhZUR5HA8GJe5nOdlwcwDXP1nA6/XMmnsaW3Z2KS3Nw2PNNcpIg76Bif2JyCbO2rEYXy5wDdvWhE//K4DzMfpqkA
WgCWiMSQ/YrlifyYMpjnsY7B4HDRp36BsfOgjMlBkbz8pCeI0TFla6QnEP3IiMonyJU8s6DH/JkUzQYL8Gj56oDvrkVaDEgB2siY6qxhMZsv65SW5km0HeuZ/T43eSQz
WW8+9436aC8EI1nKdESQPvwe/321SDd2g6wzhR36yJKaH8fd/nRwV8+P61QjuiWXFd+baqSZPUB6u07IDIkWm6X8oClxTrth3X8l5IVSCvJk5EWINBUCNlDDBZOMToVk
D8biZ95QamYHjTqmlFf7Ae+NTAbOGhyNjPCFDrKIUhWJFqbKtM6JhWSEAlUu5XGdCSE9jmII9LkFSMmlpIjGvf2aKSLvRm2EdLowZ3SwyBTEBbqMGITZpXMYdPpJUnxw
qgl0Lt1rnBf4WM5qNH5S2ZVk71bv3giK6xJiK1Z1BamoFw5vqJBtYyJb4UYp9z3zadpHr0AjFM070Chx43seh/vdwVo61jeKZBI4p6lost4En0V4wDivynwieF7xQZBu
/GHghek8L7U26vLqlIBRv0EXtC4PzaeUVxZ1KXFevBw8gm86R6MpaeKwwhBXwlCx8ONIukmpGfePWQnpdTpTyIyAYKt/EdwsRFdc4QLE7ePE05NWLjGkNd7kPAY20vaT
EvooZYnc92/eIHAkTG3/nZOuNI/vjyI6mstYICj/ob71VhDgM4LbU1HYwsZwMMR7uoTp7sGa9zopqU1Pn51rvWg5+Vdkzz7DioHCO5sk0tKZkjwmrRFIhPfw2omYox0M
DFWp1nG6H0PFocUWNtq79iBCA128iQt8P2XLk6LKLOa8JvM84bQz4NySLvPN9VJPxjxi3yR3gifOUZnjEaqqGEhJmJ5eXwKnzQ0kXpJzjMtTn7x8n8PRgHp8lSh010Yl
n61mMCloxSXtIny4cAKiUqtMNo/InK+sUGL6Tv/2Vrvy7i09Qq4reMHrI6iwT4oDYuDj5dhSVENHnTVT8/CXUAlQN/2lpUe6GSJ0kadzh4ylL+Tp7zBJR5sMeDgzueBg
BcC1XEksinneUTPeWY9M7OKWvoeXcSr37v/XzTvC6FPbW9AzLo2X2xG1i2iPLZrtS3hlE8t+uunbM3idR+9VHmfFTZLrm/PJwPKpHoBIcx/9FCm/fX2PdTQdQ4pLCau1
9ULX7izBqlCtcAqxuK5MlTmJuDhRbqM2jQOnNFT5xEqBBEy5qEWFtoVVI7Hr7z7Mvd2im59EZiX2SiceO7VD7Gi6WXcj6OyTcSXwwwdF/1DAUsA3pCbVKbW2J2fRMBfE
mVTQQ5IxCCAlLXJjw9ZAttfWQ1k1nwqRD7bUhRwFzH+SKiWQHOOd/ofagBA0/9EcTyJxRmtTD501O2QLhzi3lilMBPaX0WGZlYPUz9fOIIySKiWQHOOd/ofagBA0/9Ec
EM6cYw1unrmOLjyU3lRWlg8WxiWmBYMOlGy+gwTB5SXIRvzAhAdgRjtJeCady9dzkAzfEKSf3NEZ8MZ4ZnPk5fvdwVo61jeKZBI4p6lost51yZtiD83qVLhj8MJ0Rbit
HC0m31TuwHvXBlTCmi9coQSqlfUOvGeIkz7oTfUbX1SsknoNvn9eVCiXtBuMwXszDLbXEqjJV0zEoFTv7+ekBJct57lm+QnLzqAdSTdOEPK6+sawF07S8KmUWhvtPT/m
GZ6A76Yug2Y2WBujFVLh8TSRKG2a2ICDMwq1Lwyr0wYnA/9Hcgl8Utx0D4Y5krY0LzpU+cbZvojUcIfWr+JLtnitraPYtkzWw3tGq1DySstm8hLqvX1a6gJCGxaCf7JI
T1Hj4Yrfc9WP9OapMxOulFHgQuSzuCvfHuRDPkEjkk0X5A52/GqNJEItZIXQ0XAs+zDqL2d+8VrOHRG9YCoB5Wi6WXcj6OyTcSXwwwdF/1DAUsA3pCbVKbW2J2fRMBfE
mVTQQ5IxCCAlLXJjw9ZAttfWQ1k1nwqRD7bUhRwFzH8IxyT90WZ5rqo9wzdhBpUfBAETcqcVlXzq0XIF/VSytTcaT4VzFVg7VgTpedoiLhVISZmHkMhG44MNOBZvXZIS
WRqjgTTB3g82se8hTRZSv03froSR/mC2LENsNHvaZYGR5Q6KYR8+THQbRzHEZcbDeqAGaPgq92h8rZV2M8M64WF2V5vjHAIQrjqKqEEQD9FzQzi9Pmh3tvXHpLO0cTEn
01CQhiiPG//ZX/3ggqirHjPgVw1hbFlJqMlIZst78wDjM8plE8LeAuXHoBqzpqxUHLWAwtxvvy82rQJAEoF+yuf/AowpYykCplUpL4jQVADJU9fKX03jgafQuy+zwVXq
8A+oIJgXSyb1JNFn9/EczIfolTk7kNadx6hDybdBfqcwUbQgqCWB9RRmOAhKAxws8ti1Cm+KdmJDimJmNvIBmOzvNymKOc34QYpxdxxAAt+rEwxzATYAjpO3fNUmMuld
zU8pKatOJRPwMHUFYanHlbSQk5jLfVRqH8Dr8jnComwlgJpGd9+lm4idpMlMpTodK6K8hkyzKuT2Gzzvj/r2JYTAfvJY2zPEJFQeppYS5oWvASMfMQI5vUVvz0+Dx/hf
MLUljOg7o3zfpd5+O0yoxNtZ5RIyxAUOEE6K113JTtgnfNwmqj7vj2s0nlQTP4dALfb/2oK0RRUrF4VH/BBAXePWqdzV2mvwUWkjm7LtD2uVxJzS/TjY/sWRKmFgqfwS
M86v6EtTY3ljPYLkCNz2PSMUfUAjxsgpwadL5xJ9/qogRj0ip1GCTUMZyzXgb2n6YmJ/GbxJwpmrgL6tKQy6fLKjoCSX6cRm7K9zWoT4eDedj/G8uwaf9AOV4jQMnq0j
giR1WAppcKd6NAActf1/eD+B7PvnkptxFZ8b+Ri1+47WwCT6jy/le0GZ9jdIwAh82LHLjmjwikChatMbZodDqbewTkvrChs0eIru1gCTgoW2EA3B6kyuABEJWTC4/gLG
cQ3jFPeMldEdkFGLgZMWHmocq+KmA2hURIvsiMUQuT8Yjqh0Hgec2pIfGzphhAeDOOO6x8xr4tgruW4QtKZQiqsTDHMBNgCOk7d81SYy6V0OEitbDofc+trSVMwizKkf
U1x4+p9YuFHfYfbZY8J7Xt0J4Or494A2U4oSCGAbTg4UXgvMvaKjCnapPKCayCPYhUEOHIrn/DLdLqPvTwGd9VzW4mpQnI49nCWSZo5AlOR/NKvoeTeX1vFT06haw5J/
PmiJ66dlz80yQoT/Tje117Y8OJKVixjTVaPHUylJql3CCob+QlbDXP6frxAQKWmO0JrIvHnEXRFsYHOB78+nGxFI2qbo9EtQBrKPBNwlNdr4n7EA1dNJG4kF32XtodEx
hXNLGPX+qddl7zreoFheLkaZKsDkcKqbVWseSa4u4bxHIcOLFeeYxp2RxFkQt4JstxBk6XK1oS0j8ifoiwJEj+rFFsw3QkeQxmkmDD+9m5x+gC3ILgeVj26iQwdcCSaD
rgRxYp2cpfZS8DBuReWCGUymsfJqCl+0O+nhADGLycKOye43dLvEvlh1LWxR04TZrwEjHzECOb1Fb89Pg8f4X8pKrr3LPdT6tz8B0VrrugHDdKx/UjfR7+Uehzn9o0qi
0HsFst4j7MvNgoXKgnDLuXfpnzSgcG/KCQ4ti7d6b6N1hQa3gTF0tVSRQsoTYooVQMlBCHzRZ/l3GrzLK9E4hB0PETFlZUoNeVpImJ5gPdjQMyo9KeaK0hyiVLvYd3pr
DBK2Xv+/J306HmofHR/jAJzTbzP8mvQQzjhdyvhHBvWVv1TFD6h1ASGvY7zOhIjiELxHQEZKRsioWIpu/UfhimpYidvD0ba1po5pWrg6XDzCXM5t7DxOU8JhlLOMNhJd
q9Yx2Dn1az7L/iD5SyQp0nxcI4pq/K6OGQObcKjphmxSX8bcykQZEA2UhoS58RODMFXI+wojHZZvpzVeZ6Zqva1jj4V/V2rXWmuvxoEbxD5Ar0OmlJcNYHEevd9zvb48
dxKuGaOgv03Qcc7wbDvEzTT1xf0RGQTDx1kwYSlz/Jj+ZIlNs1R1kuBiem+oqHQuNIOC9NQU39b1aNO70XnNq97PqzxNLU/Tb1xAjmZYNBKevV+ShQ7SDjtM+0oblDY3
v942Jt90JWvqIiwQ+XvW5xEkD1qGgngpo9+SSZujQI7QsjjY671AwMsff1ThcfkdVSXBMv4+mnCNFDvGoCL5aMQsSY1qLxSA7rCnsQvGCiNx2myfwTS+ehMl0gnaVwkq
yX5ODbBAl7JHwaMVpaW/JpvyvjOnWpfvUEptvL3XxKwsjoZAaNS8iL8Wb1ZUPPZHE8Y8oQXE4qYFnPypBC/jVGxZoJQ7bmfNWbG3rvazcZhIDKykRGYmKrPPd7oOsY/E
pGDVqHv1RDuBaMHiuWoOSScwRvG/TeB+p+5vgkvXLfFMoP0YxmBLuzS3ElcEIehhMSW7xWMQFO5Ti7otKJG94ZYf50x9FHB1aTpK9yhAGL3DHdxeoKSggejdQfD+0akB
Ia2UfSKj+7899im0C6SAJuNoOJPA3VA8zIwHqhCbpxu0xghmd2IbnoWbw1YEOwOQ42g4k8DdUDzMjAeqEJunG46BEkjFi5Fh4VHp7E/f+QPjaDiTwN1QPMyMB6oQm6cb
RajST99pyQ9MRWKcejdBM1DrYXIv3C4+HjdieDVEx6p1/LvTr/DlN++yb0+pY4mCdps8ZQmz4iHDg9T0JRERdNlHSgYhaTG4/S9+QOFcNCMiJdv0prQthwBRZmyMJPa6
fQZQTDt3R4tplXntaBcywp4sSyhSvC7VWEX/g/g7fA7OQ64FnQoSgwnYwHNslcdCmCFAa5FdUQy3h7pLzkaFaOktF17TnEO+VybuVM30Cu8Sb1qaLvV4KWltnxA8sRXG
tDG/jsm2KQFM6eq1eJY6JioQvDEJB0IuYgBPAUU6YdMkzxCuwcvW/wz/XiKz/lun0fWei8G3EdT0OluRpDxC34vbKlaqbQzw9Q5+8XLBQpl8OyiM9wcgQPkhQdHBRp8N
s3RHVrEJV6JZsxxSxTxxIerFFsw3QkeQxmkmDD+9m5x+gC3ILgeVj26iQwdcCSaDrgRxYp2cpfZS8DBuReWCGXYf48SLFFMbfxbXcHKW9K8nSY2tsv5Vb4r0HFZIOMYC
wzZ/N1xIYsaNcMuAziHJ2G6GqcFsRpFfyHS9h4ewoAaxpiDIXmEccCxcRWG3vp9iwk/hwEgZ4hzenQ5uax8Zf7KjoCSX6cRm7K9zWoT4eDfhpr16kpypR5Jpm9pDH2rI
REvnUJMdF/HOpig0putXOqOb7w4Nqh52fD0RcdGMvjxAr0OmlJcNYHEevd9zvb48dxKuGaOgv03Qcc7wbDvEzTT1xf0RGQTDx1kwYSlz/JiAE0y+D6KHBFp64Kddo00h
3vQPSTuaPaRutSnNIQHGpWjkv7jcwYRqR7qyLEo0SpJbKLkdLJtf9gKzHUxX3kfju5ZSGJMI/+Bm0GrnzNQ9ZpDjfnEWZ1kiUC/5V8K6rzmCJHVYCmlwp3o0ABy1/X94
P4Hs++eSm3EVnxv5GLX7jtbAJPqPL+V7QZn2N0jACHzYscuOaPCKQKFq0xtmh0OpOUTuy9Pu3dC5tgwLqNIUms773uP+yMUB/G6+/nnLJKSPcROMust00eF6aps7uBIn
Jb/hYq1zlerW+bvxDK1Qh8YFWD1M9UQ5F1HOtiuNeZ4yv7VyDDs4mm8O+ZB2caP1QK9DppSXDWBxHr3fc72+PHcSrhmjoL9N0HHO8Gw7xM009cX9ERkEw8dZMGEpc/yY
QeUxTXicxKmotK02CqHn8N70D0k7mj2kbrUpzSEBxqXT1tye0NQT+f2UuQgMx2hSh6+ysxzn3s64f1/2Jvevs7uWUhiTCP/gZtBq58zUPWaiUuWc9RzQgrkJm/FZTHut
giR1WAppcKd6NAActf1/eD+B7PvnkptxFZ8b+Ri1+47WwCT6jy/le0GZ9jdIwAh82LHLjmjwikChatMbZodDqUv5/u7eJ/r41IZN3iNSl+GkU0Xd9WrBo15vFUOyvoO0
eDncvmPyYaj4Y+NFRXGRcd70D0k7mj2kbrUpzSEBxqX9ngC39lgfmX8wKqy6k7w1QfM8QkyBVTSoTehBbSYbLLuWUhiTCP/gZtBq58zUPWYSHtzlEgEuwtMsIG6Gsp7C
k9ynaJ8u9gVtLMlWtHiGmt4PD0mRwiU6sgQzZflO36BpvjCY/53hvG5OJosQtxfY/s10dAT+cCH9RKBBzjWRACsxvMJaSbLUP2ZoQV7W1leDX3Ziwb7zOERFaog4cVmp
Jldd5gB++6OI5SzEOKtmtGi6WXcj6OyTcSXwwwdF/1DAUsA3pCbVKbW2J2fRMBfEmVTQQ5IxCCAlLXJjw9ZAttfWQ1k1nwqRD7bUhRwFzH/O3swQjO8A1b7YpmopS14K
zkTQugw8LL4PBJdY9sFcMvx7xgKB8o2lQ+rmlUzZqQQUn06l1VV3PmgNH6TpipAxqgv6FUgs40sidC2G6uGL119c051+VHmmJTo4Eve5Y5nTvqHgVyFcRdVH2SZTU3DW
83EApTKG/gBHg9z+46rcIul6z6FmyzVb7i4D95/vz3L1qAjLo67/s3Zgecg7+SFU0WFSrp4PhKy+8hXYEvUZP2uqOkpX7ahI7Bycw6oH6EagsmH0wFY4zkpMdpPBAThf
pO4wWsgl1fiqlYMwtPqGuCfnL5lpC4OIsTJW2H/zk30l1A9NoNALkPVQUBWzRHebUCUMjGTQVTDdfrx85zadrmTzM3vy47k4Yu0UiHjEA4vPVVZz0DRn7Zu34CR3yqUV
ybfnmx3zmCCUGb5Uq4yMXny3fRikfKebptwenTlisQ/nA8BgCnTaHBMc4SDPh/6/GeWr9gjhWvpjE27hJgdZs0cfEtZkouAfhY34O/ttZk6DWiu9AS7YMpK2ZdSgIJap
MkNqmYnD9BZKwZam3w9xBKUwXcNgOTswNuhqzN+3vmK+tWtkmYPdaa0dvqjfeVAbGvWHomVA4jHbtD2IsDDS0uQAwqZ+vnWuwI5WDc4ejGju4qSk9xw7R8KycH4GuLsd
1tIh5L35srszoOUCmqgnTjVCqmszmwYJ4sTTeMcXtN1xF0bAhr+TbSXKh/2RScjLTP1DiH2xLeulagaaK1ao4RdCdRJ8Jv7HkmQwKqf+avjnOv6U8K//sfvs+tro8KFG
hON7lU5Fyqi5iQsp339XmsiVPLOgx/yZFM0GC/Bo+eptThrp325PoiG3zV+tKAeYKjY0aK4VEwmjef70Pz8nk3DtfoYr+pLHgbowHp5dPCD6EPZpLdU1odmQIul8UFAo
30Be/yMXWYTg/pDJd49goBx7dUW3CgsyO3mgI0016P5RC161g/wPnekX471w94GatVaB6bFqzPIlAHl+vWKLs1GFKo0oqAj5N1fbg23V5d8srJCQp5fESYd+W+afS9ob
D8G9vJ5G2zYxiHLq4Jzn5PBBh2yhlhmc77q+5O9g6hXwn+dKCTcFsd5fVrkvezLxNMzAUT/g6JXzKdrBt+UoKlB2K63lGZnF1lR806OVgleqIM/8mPWd6TzhYRewAXl0
oBZRjaNYkSbmpj25ND7T1Cd0/nMAG8v3UJ8Ld3vkBqzygPQI3grt/Q4fAEV9uHyg+tJHpcNldA+2RBKMRmV/s1HplQL83B9InrHvzbNW+UR+6MMhxvgFCkRWH12Vf8pE
XRSZ/Y/17mVo9yRi+YyAec54IKSECZvg+aVdBb+CQm6DHnrKyYwaPTiyT8qpt/GQNJbh0z9dTosG8scq7ABUaUz3dEXNlxkDQfYpLkro4EYt3XhM4uebSjp8xPPOb0PN
RjU/iRvXO8gBVxuJ1gvllQzHqjghXTpapMPzGvETAwYv9UknuPR5t2iTmjQKHlLmOMUCPng73wi1WQLk4VnmcsuHxnoe7WHtrcS4gtFYgP0KTqUGCcvqA4Mjs+te4Nhw
Z05+5LSUb/ypXo3weV5SunTFn/oCO6FfSaGMwA3yuNjNJwnAjJeLCq0/Old3jGlOe2B+Kfhj+Z0VBtdMqGJHDIKj6HrXl1oj/Ioq0j2DfsXSkyGosaYmo0qn3iA557G6
V8E4Frbmml6FFktL7KhvjHh4AYVX52c2JLZViZGs5+LGYLV6gEwzxfsX5LJOxWGooy//k+YjEQ6jyQjS+mnBXF4dWv5dAiiI6Fh0Cm18K2Gs+Wb+Q+JS+yF9h1aoRsdg
IfN1x7FySUZKdGGXiK7whtxajn4FTE5yLDKKrAPB488KYYoCAUx0zV2O7+27EEYYd3eSJCEGo/5w7WqLefq51n/6ZyGM3YmNwRPqnqiXX63iQq1GC3kLe6TdBcAFqqgT
7uBo9eg4O77v42x9NorWZKDOChhUPelTJmFl1JZS4CL8z0Jz7BswFciWy2qREX8dJtWdXMOgwmtV2UZS1zVJo9ELroBpyQNdfdowFQSde19sXO81XoplLRaq5UbhgmPf
Aiinncm1/KBb0KikakpHl6Ahk+8UQC/0Cu/TbuNl+p+3bcwWYvCcYzF+1alcWyQEWmM2QpTo1oLiTfvfflOwNBlsbd4dF5pPhUhom6334sMigKMlg5qJy/20yKFO13Yy
KhEoGjx7fQqKawhKOROjwYiEZWdx7xIfUZqUMWZMzDqUVKY3dyIrzBRcVd7tiBUqX/BUeaXwwjQ7bteviPjHrc43Rdl+MHE2TknsSCiHAfr9V5HRWYopVFDAjYkwdXNF
n1RQgQyquzYuhlwmPD2IVqiO1mUkpoPbcfg1ZgK+1eLfCsuqJRNtTp4AFYgnFZHNmAyXTEStYCwn9Xnr5D7dkitMqgt3eFXe/7vKnulS0igm9pcQBmePGBZe1DZH1UPn
QxCc6A+4Qz99jtyrMjFqMwmZqTzbAh9TrgOcrQqgMXxromQe106pb+zladtsAITHvn7cVLSLOdYeHdvt7y3nIlpgZBaB/h25AaWZHm//3lQP5TxWxq6ddw7Em5AfK1Cw
P0g5re+TdPUlthK0bjYdCz7zBhnrTNVBF5YCO6o5AkxC2wJKp98HsbKOy0+wAWHI4vL2A38Ea1n++aNkfvVo2jt22lZp2EjHvkpk7WqFx9KbwimK+4dIsrNySOdOTZft
4vL2A38Ea1n++aNkfvVo2hTEwXhg826fhD9O7cedgXcBfFH5JO5w52EMIq5N2RiQRZiYRnvluPIhjAZ5nlU7DtiUHi+y2hJEUrLBB4J+ap7uImdpq+VdpXqMvp1URiUA
OdYoXOiTIRt/Xi4KpH+p1khWbp5HpUfQRiuMcfzdb8F7iHvl0zp2WnP9/VWxwEfAw6gF2MxeRv19bbgpSJwQq5b1vMuCqpWK1IQIFVP1X6xm8fQ23xw0uynHtbQxKCPi
TqHXlCmGoAY74h/oX/jfqiIkdslwyU1QMLDaR5vFrl/YseVnkuUzSFCzKKCiMhffdAYKVPekkVBChV/Ib0Boy/tuP5YPHjYRfz/759xNxaEywQPyA3Q1ADksn9sBEwXp
hNJgPNHAqPe23AH50LNHfx/nO9PlC6U2ArsHNXQwLzpl+bGdZV9zf6Ea9WnlGZH0UP1XLIbqnS1xhjmEHwhYOQVxyUFA1vA4BU9vxx4ADradwbiLxp6EHc8aaFoHNFfK
bA1vchbVQ4kC0DAi14XL6pnEnT0ARfHTXTcUs9gBjLOq2ApubPqutKjevsR0qq1+H0ERI2CM5t7tkKEtqvejsspRV0XsRq8gE2MpyVHeske1xLLKJFbCgUXp2GxSH8W/
tyZwwYpyr5V0WbU6ZSYVu3IAQKUJhVGuX7ZO5/xSm8Ireg7qbuZ68sMMQ4saebI4GoyhnViazPdD+p3Hg8/2quC697PosMutyoasbFzXTFVP9u54EfayCLhMIghZXsRf
DI3cKhONt77+zm1OzvRaPRicNgYTl8B5WRP1qdg8/pVkfwO9XhG5xQp/77lEVl30o9DDHsK7wJwsSGQtUXym/6pWGHOS/Uk4kKkiPNrCg6PCJN1+xcKo5o3/fEvzFxwo
BCu6jkgWSowNu+YBPmMIXpXM65Ppp0BLeS2QBdb2IAWabB3NZAB11hABdopWeExtTY1GZLxJtndBnzp+Z8yLFNSNxBfVe06NOhSKtQ0vQlt9v/0roSEoTNXgyCtu0s9z
j/+VgbAXVS8My8lc3OFAqgBzVJHNzhptf459CDafCM3MXHAIqQ9gq5MZE1rNCpawT+vPbd/VyF5J5uecUFZ+78vRBCCOXugEik3HQejdzdA6hl488YnM8GbRH5zgOAW1
dTFZ6iCYsExm/rH1N4r5t1qPRRVXuq78uYQrQ70u3Unguvez6LDLrcqGrGxc10xV/Mp+inORd8aKVxwzxZpXFU2858IVh3VYKTb7uRDBdtnHbSSKXfpk2iraxZUEDFjc
iDIfPHup8nqvpuOl11FGPEAhG6bC2/pfSDoVFcfLXzX7bgm5K1FxyXcDeQ3MokARrLSJts9wnTVlhn1GlNu+VDHdCHZprhqUcabl8fpRQQ3wBPrdCsNisyMOwbgnM55X
KxphWoFnXwa3AB0j13J48ylNv6sxuhMqsiCfWrH8P299v/0roSEoTNXgyCtu0s9zj/+VgbAXVS8My8lc3OFAqgBzVJHNzhptf459CDafCM2j3JKdblQ4oeaaa03bFI9o
3f3z1a11w9kg2x58/pkDZMtzPR7Nc7FtSWw2HMfrI5+VxJzS/TjY/sWRKmFgqfwSM86v6EtTY3ljPYLkCNz2PSMUfUAjxsgpwadL5xJ9/qogRj0ip1GCTUMZyzXgb2n6
YmJ/GbxJwpmrgL6tKQy6fOq1mhtiJoIJk7aKR34xBGQDm7lLzUplA0rA44bAiry6kMN12X4y+WHJLGYvqYDkpjMNXLVJ/IJTwfN3ejiGTdb4Mq1hDvmDnq4FecW2Lk9f
U1I5hFlsrd0WbR918dRLRJeaOQXBkvC6BDOfUwJWoXVHDV7861RdHN9J8yf6ssIWVEeRwPBiXuZznZcHMA1z9R53WUhuw3LbYQh4KutGdE84VRCrZWhcdX8ES/m6j9zZ
6lWy/MZ4F5x9eN6muil42RwpKDkOmj61EnKrTH5+n96GM1x2N6aU9T0PmJHCGgFU6piYt0U+sJJB3UN3mfk4REN+v3ygWyxZRL2KKf5q2dOxvDZbWP+lUPnnVsQBK76W
lk1wvh/RY08FhfPFze0y5sUL52p16hRbNiZxqbXUY1ah2M/dq1A4j1p7N3QjZybGQ9WkbIFFVhD+ToSriehvU/dyYSJ4qYRhSd4sqtse/qBjSUoqNagWlUoBRfFMIU3B
4K/Ayx6vC/IOVWE4oKGYSIT9Op5SRuTNrtEDR/hFblqskYNY5ABeWZXiuDjDA/ajHD3VCM+gI5J9wWr+uAaxTCxH2zNgV7hl20zpzOZIvnD3jmLNfIJRPZCrauNDvnrc
Y7GaUY0zSM7Q/ahM5YDsOSJ6teLTBfBM3UQk98EyE4B0goHXblBakMmlF3xAH3xdIEY9IqdRgk1DGcs14G9p+sCyZgH/Hn3awrxEkaDWPhVmsOfDe+cTRdiY6Oi4tPke
yyFiB9K66yhHpA+CCpio/3MI96feBnKaCJUtuxzVOrYydSFsHv+n/4T1Bg8m2r5KiQkwG/7G2spX8Ahzu2tVPgXAtVxJLIp53lEz3lmPTOzilr6Hl3Eq9+7/1807wuhT
21vQMy6Nl9sRtYtojy2a7Ut4ZRPLfrrp2zN4nUfvVR7cUC4o6JzlfxK2ZvVZPw818PRlqdFb/30uUZQO1egKNBDkW2vr4lYOQkdZNZ+GDI7dtLINd4DMYlKR1BDZSaGf
pWGpcB9+4nvAp4Lp3iHTepe1fvKd6KZYC7TwF0yiVOgiDnoMfjyRNd713wgbQSSgfMhGgytLRR7EsIbATo17qz30O1phkxycJFZoIZbYqwQXEwDbdZ/KnLdRTWNgKfio
4K/Ayx6vC/IOVWE4oKGYSD5RPOIBSHIpdGRR0T1L5vnccFftsEsp1ujyRZ3QxjkYoPdZ8/N7Z7YqOQFp/xE/Gvecroq90yIw9zAHRksyw8s2tsrT9LLo5Be1BKrZHJR9
Hk2mjL24S19KcqpZnrPLvtR+tHsCe/bgwzx9EuYrN5gaJrqhuFmMzomp1kzHfUsYWPtetglEj7TVwFF6VAqXaQTgXDNFuj941W/j1eUkurlc7oWW7Y/y8ffiplxZ8gui
Z+FCvFp/9M49ynNbj1RaTmmSRyme9F0YwB3caDk4D/zIIUDa7hNstwYmg3W2D91ybwZQwOu8ZRmvecUEA3dkxsiVPLOgx/yZFM0GC/Bo+eqA765FWgxIAdrImOqsYTGb
L+uUluZJtB3rmf0+N3kkM1lvPveN+mgvBCNZynREkD5MZYZ9Nq4NxlWKSIsfuZRmipXSRLC3M9g90lWg/n0ED/x1mjbL53e4T+k2Ni0TuSc1yN+3AFHc7GDYT8DywYft
Esfm29ISuhkHKwzr2qBD2h7E2SEE5gkUp7PPrW9V81AYn6yBmD5QANABpfDDUa7y+msowlCHhtO5vZc3OVWFf9fRsDsxsrRobRul2lBKeu2fDHtpn+L4yLvfEz0vhvhy
+2jbN3KV3GoGausrhIXwFSEvudk7dLYD7qU4w1V+LkcQEC3m1nkbufs6dKeiCS2VIAMJWUev3FlIjoNgvTILxqV1lWdSDf83Q9XBa0YUYv386bQ1tNgCbQov7DRIq9AY
YGENO+xFa3GpEIkf24FQXD55pTFopZLiFsMmzgZABnEswXMI7f2O9firRTisXmmpg029Rhwd+8pX98oKzM6ExADvvtNtduYLVUPyDwldiolHOztmUqt77Y8vRQz3DqR6
CDoKqkJzjuG4Zu7frBcXItu5IkXCCzq4vEAvTgg2Q+MyxpA2tBYaCKQOgURO3CfljO5x+zTRMcn3t7wxDbVLiX4AZrRrR0oVIPXm7Hk1alMn0w5gnGr4a5Y/IAEhoP+5
L3JW/SvX+5iYXkXdB/W+8Zwy7R+5U/c+QadD+da7BqyCl6Df80HXp3JLy/vi3IKP+hD2aS3VNaHZkCLpfFBQKE6MBQassDYU2z/gLQybvM0NQLygcwA8J5O8HAnjnWvl
p5cofhN8C1K6jiAKmTsNhasA9ACf65dIZacfsQOX9IAu/Tlu2e2XhEot15cpVkfQNnoGc4zEfF+SofxrrYF5GUKDj1uP3by2oFGuvZv15R2LvxeDWT0xL/ed9QWPNg/U
Z7MXkpVJ0EyA3OIHcgC210jVlZMytr26nRLGXL7gNB/bYPWoLBflH5po+OH9UoaV+gfTFCR2OmkTn2xLOl7y+bItqFne5GJdfj0Eu7rejhG4hMsy3C6O7UReWsRjPZoK
RjU/iRvXO8gBVxuJ1gvllTcq2n08crTmqUieq4JFRBGJpSzQpda1/gF3NH7Pg1PErDh2u0IKMTAiEfDCuCx/UR3ZVk6zNTcQoc0dEha7bzKKG6m/Gm5ZSJ7/AKR44TWv
zrR3BCUg+XYZpsAUs74ANmFD2xpSavtBikIPm+VcIR2RKtzMpSn8r69URwMM99JnbBTNlM3IRIuEiSFK9Um2kvEIkhr7bEkjEFdZbU+KCw92SEuI+veKRmgFx+e7HEMZ
J4Yl08wJCDUtMoXqnHl9roETXsM9oXDSPI2YMiwEMA3zdG4wp5p8saElvN2/kW+rHwiPODcvVmQLfUDVcH0hDaNPQ6rgg9B/Xdto3IK1B+DuYcHnjlxOy9rIlmxYvM9z
9axyHkJDgR9QfL2yPiG4lgF1ujq17y08AffFzLuIGzWA0GMAFpTGlrgpQU3uNNd/Olb/5eQAICWCyS9TIhTLf7uUMvZ8B6GyUMAeLteosr1Fmoch9+yBLSbiqzaIZZUU
3T6L+AtXDJ63k1P/kC5bsYeelccWZaZXulwBetB9iqqc9LvCFf+Rf2TgLe78JNf8ib+8ojnw94BtJmI4+zYGqpu7Hg6T6AFgKgnwmuKhwBsNOdObhqsjZThhVoMSwQ7U
pnwKEyHaHHlsfGzFda7XvZxsp7E1/Sz6qQbRd8lYxFK+gxw2bl+jcIDkEW1yJbzbBhdQgNalGVDIcjZ9UK7rEsMe93XrbqWREKwcOf3FDr8q+5XPyVeeLVnnW7h679I/
vLq+Q9opSkDIG0HJ8vi2rsyhiiPomifOgP7oNfyaZeRvnPTxXb2AeD/cs944h/NEXve3ZP4UBuiRi3w884LNkcqGHaCnUQ1BNJSevaFL8dzEeS5Zj/8usOfFGESJzl3h
pu/s5OAStXkuN51JlPubTk+URLUlrG3kgRH0fJ/1/2yqCG508idA1JTArCf3I8k/VLi9cCfMOOcUVLekzRtf/G6iRcsQA7dhK+FAw5ughzBUtLnctlMZdZ5wjqULUM9J
kXUUVqlAWia2vPD1WFyJnhbITflOH1QlCz3MEhA5SqNFJ/23DaAn69RNX1Nk6mfwUeQZbj01Z8B9IgmhQjgsmB5XFj9jBlBBFxe1C6Z4+1wEnVTfqPJxh09B7UC5hDqp
zfaiWH6wiPp+XfP2AZDwPxRvkkBYiWa+kjoVmcFepgJB6nQVU/57DEFTCkjLZ6swvConluK+B+mHXhwqgfseJtJWDMWt+Ubf2U7SFshDvQK4cIFt00qo2pggxTvQXAKU
UawvXzau3izMxjLnWrg9GYYxaRvxMtzSM8TRfFCj+/oLzHMysCcOqWi4yzrXyJRlbbXeyTcwql3wlVa8EM5KgY2MJ1ZCAmdYmuIUqsAC+nwhRTl5j745xzynzVobme2D
DoFylGOaM/l4jP3KnLH1D4DLgxVFuN3YxA4zgpc1s/4pyx+uH07S2KfZI85QcQFrqNiRJ/Hos/mv2kuiIXlCiAoGfLxnF+lvsgfuoLX60LWgUTYRb8cWY2MSMiYdIUXG
rhNVQ0I6CXcDULiXgJNPoEwq0WpRSz0tYn4nycYPj16d7gyfRw3ogY2nRH85LMxm11Y6e6rkyhuiTTsQSLRVOr8+e0wvdDdRZJHagGu2IWYWvxJIWbc3ZHKHozxId541
USOPcV3rJhu9fmYgXcNimiluh2Ft4ZFEofjbUm8FbksJN4jP8qNm4yAPMtlllJLkBAwY6RZN6jmdX1MTUxmPPe5BUaFwC4LaZXA+Z4pWmRce3PCipJS/Tyw8kr7D5ESX
4ttRz/JXm4OoG5jis7hKafvAtkejPXT9ZfovzIxt6olSMEDMNn5WzS83Lo6msNw3YRhrKHtYl64hm6vCGN/IE97lsJzJVFgI1bcyO7BKUxsdieDYzzEjw4hDK3hxO7wn
YhSGaVhzlZKIjjuv6NN2m1i5VPexAtLYOG7gQJ7HjrTwxXVVdtUtGP+hBIgHbuGaT79xpNYCyE3CseXmHQV7Cq8mqJWrvlD25XG/oJMfJx6S6ko2/djHT20omYPIvnkG
gW6ql15TdEvv31QAft1kajuLbEqByNu03GpHD29iPHeTvEXDnKqSjvUCZ6wfibwpvayGE650waITGCvNyWPhcHzuaXVgyI6QPxcizTYfRLqhxzCCRAQoF4XGuObqjiG7
s3mtzaMtu4aLQ8f/1oRJKfcA5QW7i8RHIwU2yf9Eh6RdobGWLe1AoT8712o5fjCdZORFiDQVAjZQwwWTjE6FZNk84A0Clgj6mUm2Zxb4obQk3Lm4O8tfX33qNQVwdG6p
Lr1jWZywBnEvPgijmSz213o8TgEYB2cR9fuplOtxr8Z2SCch26hrwKXjmuJs3NeaC8S8DahJeFBH2PjWAtu+hSJF6MJYXRllFSns1pLWU4xsCUy6yIUvyFKrXa4yrS57
YDZKZIOYYhnl6jFhLDyIKQ8gDSj+xRfIYs9SbkH93CXjnwxNnqqZ9VgUvh1/crtyyVtDhr1U9h+W5vsayz6MgSQT3g3Xt6RbYao8S3nPdviP1J5V4kmDD06YvX7z1/Bo
xVxaMXLJDHyAQFcrLfJDemOrpgB2E3mPadGWNcNY8jWzPATPKNkDxVsvp/7Bu6BdFHRf6vhldLLSbRdlYlWYwOR9M6grx736UQG2BewKfGVS2VR9a0q50+w1SgFBdVzN
gGfHs+nd3hOtyeAg5itXi4j56XJZ3TMAkZh06wauBM4J7Ap+TytnIxRfst2vwF2Uv5HeK2wSOAxINmyqBSod0Wry4tk1qdpGuY+o4cQUZXANdxCEic8CAhJutS0I9FZG
8EnBATXuxs+P+88gG51sicfZSxkaBOqbLreUBg3W3+1uQbPjYaLHDYzxE7ATacLhh/VFrVL8B3MXhLLOhqD0/4jP43MCOCX6GDFBucfwx1SSi+QeOVBHSk19+FmMX2ix
hHudup8UQ0gHx2GKi4cVItrNUHiTRd8ith4rsMsT7fNH/t8TQpZZ48dF1dwnyXFOAvvn//YbLG+xy7LKJhlLhS+8NCB3IQaF7FmYIqFDsT7EyvkN/CIQLvYVlxTW2aXJ
yejFF429ofIDuBHuI4kJX4lOaoZbnUSix9pNywe6wn55iHKQJBYRazsFHAslmHosoPwndD4Kzm0jvBShSM8HxLkHH9sP5RJ9HN6qkuFV6NMO2Q893BL8vlCOdNz9BlrR
P4Cs9oRdn0A23xeeW94jDnXmPZavnoMm7e8KTEidLRD+4UGA4Ve6E3sRU+ENdQrTfb/9K6EhKEzV4MgrbtLPc7lMIk8ksS/B5bPGz6MuEL8GQzQ1E9rCgqaacYpYbK6K
N14bVA5Z9AV2V5rS7Qt0zO7qrGUoQRhESb4FKLbyPcnUfrR7Anv24MM8fRLmKzeYGia6obhZjM6JqdZMx31LGFj7XrYJRI+01cBRelQKl2kE4FwzRbo/eNVv49XlJLq5
XO6Flu2P8vH34qZcWfILomfhQrxaf/TOPcpzW49UWk4rfC9MpARL9IUJiZe5cnC2aNsBp/OJIod56RCtwr7SmZ+u3MGnVoiASZmJEkkLFPMTwvSaseJ23MULniBAj28k
rlUgAjXAB2rWHa1TRwHjF7xnvF0Z+962XnPG6QhcgwJ164YQ4AkAY7tweHVF7Uj1tcSyyiRWwoFF6dhsUh/Fv0lvxkHJ3ogpDAomrQa8tbupYMYJL/iyE0WBOZa+6UW4
XGBl67TpcTXUfFza31vFFXKbJyMnbBQxGG1ISXNWmc2CJHVYCmlwp3o0ABy1/X94P4Hs++eSm3EVnxv5GLX7jtbAJPqPL+V7QZn2N0jACHzYscuOaPCKQKFq0xtmh0Op
++QgV2gKj9yTzVY8le60AkJvfXj85aUzFJXpUqHad9NqYziiNBnNtk9U8hLlH+2DpJvhKc7dJfH8Zq5+iSSmLehpqWLqGoK6tRaMLupMQbf+ptYHZ2hJASQPwBRYtSmU
eRCkzNgzZ/OHUz6h1j3vHVj6HGBYqhC9LO5ZgmJZ+frKmji7FPEsJYJGW1gkMglOErc9hKDu4JKoJ4F+IWUlFWi6WXcj6OyTcSXwwwdF/1DAUsA3pCbVKbW2J2fRMBfE
mVTQQ5IxCCAlLXJjw9ZAttfWQ1k1nwqRD7bUhRwFzH9olQolaRkGuNA5mBmFGEgXlC8zVmZ/vVsj4ogBjskKu4aCBNU8xPG7LzH8nS8m5zCYTWdsEq1BHUluuT3zwHo6
pJvhKc7dJfH8Zq5+iSSmLZKSKOr0kfRxUpkM8A7qo4JNLVbCxAeph3y1HKprevlZz5nFCYUq+QWcn9I92n0OzZzfByAng9FjdLlSjhQUBpfMlRcFfuDpnailI9B7yw91
GfDIXuOKEE3PqnTW7X/uHJeaOQXBkvC6BDOfUwJWoXVHDV7861RdHN9J8yf6ssIWVEeRwPBiXuZznZcHMA1z9QzPEQ+FscTmgM1kzL6sEzrDWQ8JRoaOVgkX3MUQcpSQ
SjCIN0SOZrQD165Ela6knMWaWiHYxUaZ3Ry0wf+yXcmnOIRz18ZtIxIBv+9Kt12UqmiBBZHnNuYrF2dkkZinlGMI4USMC4UDgB3D1WGSyIjjnwxNnqqZ9VgUvh1/crty
e5qzhoXGetAMQZtxofcNPIcWJ1iCj41IElCq2lhHn1Yeil/+mu4TiOBWq1mY7ymwcwposFG6ze6avhNEi1Lp+ufMMXVisgPrUgSkqxJOykkPISkJP8dZR6fwDt1S+Zkt
0aV+Iw8R2ytgYjn/qFeAzXjzBGR34tJ3liERgM9HwhYeLUd/aQdRybZ5tBwF6oc+ACc+ve8i1xEiQwY4ZOhSShF7Lfkl7NQ+VVIu1K7G3kdUOTKjFCSlFJ4hef+HxeCC
C9FK3M0XEnRCsM1O0nk7buOfDE2eqpn1WBS+HX9yu3JuHK/seMPyOimMom6Ni15mNZcyMXrP1pwE3dB5YGEichw91QjPoCOSfcFq/rgGsUw0L1zLiqWnrLhShJgthLOF
1lbB9aInCcyzjbiXBCWl6uk2+56A2DG9YKWL4d/czpaGME/18SsUKGqX/yxtISFtxM0yQpxuyiTNkQCnvAV1cyZ8aRxuB/Dsg0gbmta04cX+/H8kxBfybmV9RMxSWzeI
/F43+CGkkQVGCZ/QZOxutMXPUByRIR7LHAJx4Pby4R6Bu3COp2nY9xqB6YdQQ1dbtSI5sHVuHyYKZOuMhuMDPWnovo+G+m5Qc3HRLhzn6V2L24LSwxuWZgDb1+mFcJq5
yJU8s6DH/JkUzQYL8Gj56oDvrkVaDEgB2siY6qxhMZsv65SW5km0HeuZ/T43eSQzWW8+9436aC8EI1nKdESQPm8hwE22e3zX9isOsFni6OzU7CxB/77D5bxsSlqzjUjy
7M/XGlpHhbtSMIBddf82uO2ONyzpr41x+VcT0nTr+osXloDThzwa/TVEb/lX3c6yvaYIp62UvFHvqtg0yWiZEH+ScHaiEL//gAd+Mq+ag8CSWAu39vdFiKtYmdja0Y3l
PEKMLIPx/3MJB9ojFP6Saa+GMUeWJiISa2QuIaVRBJiXpIBYgKK+al2eTlyQfECh5wk2WdB3gEXmmGDMJ6BX/FPG8GiWab5uuCYb/msd31W9O5JfBRAknt2acONvqiuW
9ccUXQWlUS2DwIJNi6zvU+OfDE2eqpn1WBS+HX9yu3KUh1TCCTVGCek5ymbXjHjPXrlAaQHBaGfgq3Ji+GDPWcCstTCup8RqzxdJASsfB018s9f+pNhEWtli/LzgxCU6
G/DRapEOhMtx4ZW/Kb0NPJ3ZHDZgWIrs481Tjc7DyJ57SgaVOXceLxXN2njaOG1nkqOa4VbOYD7MrOOSSiMnCVGPzAnX2gBNnVs21gUQAsA1tk6McgTKC2VHh9uW+gY9
U8UiKdtAfu3YRYWBoGiCeyxbiRQO2kY+YFCggo5HNMZLsXFXcd5lwSn2LeMxY99sUbFdGdvPRpPbMhfOiIOYyyOxlpvvEKHV2oJxUoDhYDYsW4kUDtpGPmBQoIKORzTG
x/YF2406u9HIWj6lmHaF/FmUS9rRwhEVVdU5kq4JMIc5S0H4qJ0HJZt4aHKeyppAJKSIscbl865z3eQlZapsHr4oASLovXDX4pX2rYqv5MnAjBIZwuTQYrJs34s2KPJF
3tJwo7y2TRYX41rAeQSW3o92vuScdnDdyULtu6ih6GRPb7ITxUeAkIDB3fOdfieKBiIzZCxvddR6ZhW1zKLdrT+8FwhHRqyK37kS0YHm8bKeVccWHhj3mIYBTQrDfPck
o0O9pQzadFIZ+A832HvNg+P7XmpDw9Aja+4Znf0y4XupaMWtKRspa24XOAuPWXeqouvxQyXz6GYPdPnzZqYOUMdtJIpd+mTaKtrFlQQMWNyIMh88e6nyeq+m46XXUUY8
QCEbpsLb+l9IOhUVx8tfNR+6Z8YAWKAIqFGo42fGrU+arOoq+L0hoKasjYJwKSbEN55yRP799ZxM9awXq9XwmoHUWXI2ljhub8A7aAvX48F7hDWled0ECgVVYJpFnXcO
/g4MpKl6G80Fg4Mk6fHl2YIkdVgKaXCnejQAHLX9f3g/gez755KbcRWfG/kYtfuO1sAk+o8v5XtBmfY3SMAIfNixy45o8IpAoWrTG2aHQ6lk0psNt1sUv6btEMtSgSKY
EUU3veUurBA8xOaYeDqkTIDq+CcnKrupEQpOEOhSx2KwFy5obFk705WM+x5gw37EwEJow4XuEn4zIlS7hkPEN2UuZxAuY/BZNVt6bDHwJoCD1cndIDC1Li1cRlfna77/
TC2Si+Y0gB42I4vWEvcUKoFshwdqV0jTkllfzspx6RnQpvDFCOYbkQb5JpytySILD0i+g+ngzymMY5PPQ+rZtXXib4eDbbvRk/WqluWjBNxZbOk3HH1jYwOly4MgECDh
1I1zQ2rmMbEwyxSqpDDAm2LwgFGk1Y8K0GWinXb+vK3gXt9VB0SEpKxiEWI6aL4taBtt0bRzvYTxhOUFNyJRwZg4H9NL9TTIriLm3DebsI24iPZ8jbV28gUZgKVmuexy
lBTRCNQrq3eTQTn8WoWuqvBklf7eJGVrh1Z55YTn3gCDTb1GHB37ylf3ygrMzoTEgVHKW0N+k52cHGWu1F/pzezWUrXEusvPOSpybARy2pI3tn99CF/eorEq96mqFUHv
NMkjeH78FQmIlPskVY2XCBs/N2RoT89Q3RmYU5E+MDdDgdN1743kEBSOdJuUDDsQ6sUWzDdCR5DGaSYMP72bnH6ALcguB5WPbqJDB1wJJoOuBHFinZyl9lLwMG5F5YIZ
bSf1HDoAdkya0HaN52DDBSqi0lYf2x5KvK+yWlnZXCj5BZvO3a7BVqF4hMrPWheNLkkgzIlTxUHDCRlWbMnDhlCUofMYW5xiWfqHxNl5SI2Dlk6J5MtVU1XV61kfdTXk
m/+8SzIj+1vdnsAtFmTUhf45jOoEBMnzdrUziLxRtIAIDOxAoa1my5zTpfdH8+U7sb/0TsThTzNndPbcDSCHpcNXkSLYzPFMLmmphhZ2Qk20Y8HK7Vw17Vg4tr1g2921
SZXdRwN4saED/s81w/rdTCmDeTq75qcLQyWkN0vgND44AdYAtOWhQHGe+y7dPVHihSqbx+omoK+BwSa0kDGhL+YNzVcdWuPdyxsiimIcC5AL7asmsobBP+cm6jO2FXTS
1fZNCT57uz4YVfWOHydrd8qIJtEmvYeBjKtfeWMCbYgf2Fh0kCJALQ+gfS+W/Lh+RGcA29HTzyHcjHXAc5UZ6mrfEDbnHfH6nK7zyIl8qYUIfKInbF1hizbQmnWRPlEX
dYyCzUbxZGlwSPrY1fLKy+G3n0x5XjPvM5gfXTyd3kXKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYhLXpyWdCm+Bkx/7/krtKE7
vFBert9E9Lzw/A3KuFaACheVu8Trf38dJbwKwOZTtAG8UF6u30T0vPD8Dcq4VoAK0LFarzn8S/QAzaJIAPv+t5xkdG8ZLNU9z3uYCpsSp9aoXFqAvavyRGvbLC44etw4
3gRHoQ0bubQUMPVuAEVMOg9xmipgVxkC5LuDEUkPLXAvW5jfQESwU/QjmSzI3t9cl5o5BcGS8LoEM59TAlahdUcNXvzrVF0c30nzJ/qywhZUR5HA8GJe5nOdlwcwDXP1
vqh+a4j6hpNicVx5Ti0s46Sb4SnO3SXx/Gaufokkpi2XarCqecCEH1H7ZVSmxRLids4GpdiN/aC618jCuv0ZV1ytit8MyIAFRHvnLIzCVhZ3dyHmb3mKIi5E9AbbyOfn
UOthci/cLj4eN2J4NUTHqt0NkXPAZ4Ps1OA7daBmsCSliDodLzBE5uNa3fJeaXqSNH9IwBj3DFbVuJWcYLCQXI3RcGMVK/AuHsHCmGxYyTyqMuTXxsG9MheDhTTpZNes
L5cmIODsZcaPuISxMcGpX/BdmTlfG74AmZVSDbzZmStYdN0uyNMg9Hwj4xfrkkojzTKcvJ+XLkQh0vAPhjIjft70D0k7mj2kbrUpzSEBxqX/GN4hz6qGij+NV0gglo6Q
N9gvr64MGf+v+jeaHhM5X4JDJPo/JnLIiQtMlxGRNb3TxNcJeB43gY+WIiSR6+XnGTuDY2WVtwdpeoxjjVNpm/hPsJcP1Bk2y9cKmC8lJJaCMYTmsDq1P3BAtAExuFv3
I9mAz3TcOxCpwEpUEuQRJ7wpCfveNZ5FQCqQODouKPDzWWalO7WCCrUhl7a+l5mV076h4FchXEXVR9kmU1Nw1vNxAKUyhv4AR4Pc/uOq3CLpes+hZss1W+4uA/ef789y
9agIy6Ou/7N2YHnIO/khVNFhUq6eD4SsvvIV2BL1GT9rqjpKV+2oSOwcnMOqB+hGoLJh9MBWOM5KTHaTwQE4X6TuMFrIJdX4qpWDMLT6hrgn5y+ZaQuDiLEyVth/85N9
f/SV4g8J5o3gcXPXhbUY7lyitNTy5+ZWuvoFJzdvIXSrE15rK/Aui1ReuyCmRJERhzV9BBu5VhiqqtRtruI6d8FgZzNBY3p5dNbhutIelQ5/9pPH4QbYGYZQiVNXYPu3
a/Ed/3NOmTUVBkEz5PDLEdj1QZ6OlcHJWnnFTrpixsUUZKPEeoCC0Hf7B+1OMXA98XVCev2lzqbym7kEm/S10AEVRkojBdAct80X6EjzFoH9WG7Kg668iMdtKXE+NO3j
bFzvNV6KZS0WquVG4YJj35V0Z/XQw58KHDzyNmrgh4N6Ka3WTFXhEue5Duhk9ljYhn5jzEZHI+KUbUQWcNNZkt9jSfrVPAJG3J/yrAdVWO7183Vf7WuULCkMOBibPHAf
VzdFg5g7t+hLyKsLi4tZYsHmiOnY8TzBZTA1mtyzRTigvqaTB+ChKogLcnHYyPA7HsrAj1dbIH3Kc932TIBksfbqfUW1OfFJq7jo35QqEKjAo6xxMPVPUWOUbqRv6EVB
yoYdoKdRDUE0lJ69oUvx3MR5LlmP/y6w58UYRInOXeFbWkNEhj9MqydPAQK+wYGU/KFzENl9tiRY9amrNl2sNlZcmtfCjcMiovSW6UvqnfwGhWeYJjifIp2Q9uEvFWaD
d4r1TYhZOC3x+EZqh1/aems2/iC3p+MUE5z4Gv52uTC5Fq3mKhd62hpdeagCJftr3wrLqiUTbU6eABWIJxWRzZ3kkJqx3jSco5aA27/9P8kDJVdsgrbWNK/sKTDN9NBe
q4WR9/0BPYVY6mkvIrTCkgDeN4B8eghm87tDUVj5NwhZA7a394F/8JMU60txuKlhYxJHKFkj7kVQadpujbfRX7WeVBZSPLpM4bhizw9kIvUYtEqvdQazTHNlULStOz5+
CeW30m3fjy51HcqaObFAhFI//+pnobNWw8BIA9ERmITJfQB+zttNneicx1ojUDB2NUfpDOrKuK7Jf7kDTL8/7TN+09R8c2zvBAZOq84i6op2d6KSA1MHJRrCDsoZBRtU
Cnjq2DRxMVwMIJHCiuzFObUeuNqhqkka99jQvPIGbXQ1xY8WCTHhz6BguigBpHPuPtTo5uDtCeU8jH+DDrpGISE9UqVocGN51gtc3DK4nar+JE108n8XqB5YVVu6Ji4t
9PX4fFhQSBZnYp5dcPLSYJ+80OvGtnT32RCL4lA44KLpFlfohYFRMQUMm7YyLVv6NsxjWJ43JvNN1pK1NcfXdDHyXQ34svXsI0/0us2bAFSbZuEofIeDz+lRaqRm4toL
eNBH3Y63xRg31ejA23MFJJXhuZqqgI9j33vKQayw9QB0jhcULdMyWvA8SyXrMEBED70c4o5yq+ZDJiDohBI5w965/mVVwxd86cuwj58DtDNCjjBbdaOkq2q6aVMh47xd
GiIqAUbgZnEWQDKeh2tlwF+dHoPSgcHsyh7GxnAasXh9ely+YLfZyYoDmhdNIrAkHSMdrocKg2LYyg7vIdwGbtP865u4ywfvvNhm3Cv6z7MztjnPDziWC5IkVPHI4ZCk
NOOYofRotzpgajA1DEag6lcei53flIGGShu1xm6LO4OUZZO0NHc6O5ouVlvMSUqx8mZvdn6a0GqFOE0VU1SaxF+u8/W18gZuq2Aqgkw6n6EKJwzp5dxXHx0uoD3bvZ9Z
F1Fc6BvRSPKSF+u/CyLTgH16XL5gt9nJigOaF00isCSEZCcrV03aziL4hFR2Jy2HGLlzCslvtjz+PC0qcSRT0S4vmxNB6NN8dxoDSD0b8dynFJaqIojeQADYQvLaZnuU
wa7koKjTB6g37mbhnWtfcltuBd/bfxbivwAtCP2z/FXlZ1hSfzlOavfEW34h9ZWpff6N3i+H471wqVpe+YmsqqnJr8k7iwp2g4ohfooeEJZmOtD3nLyHYV67axCBmaJo
DRAEO+ZZ5B8FZDtMoMqwAVSyKXBf1wxR35NMyGCIuZKII1m7jZ3TkmjCXh3tNrcIxq6oSFct3Ke1giF0tMdekgFA9YVe9s8hyg5j2B2MKuOEFHQ/fnfhD6FtyzMVxzQ9
5npFEQrkz6e+5w8lCH7ewuQdDyiLppl4UjEmwnwtXHzgkfBu9yoZ7TQLQIgTo+r4b7SCGpH+yVqW41ov/fidNogjWbuNndOSaMJeHe02twhRKGXzNrtA7dC2sc9hJPE6
AUD1hV72zyHKDmPYHYwq4/s+UeeDfO7BQBdYB+RI1cPmekURCuTPp77nDyUIft7CFCRWKT+nQgXPaDBmrGli5CRVCbtj96897DHUuLeCuhFNtERRuJD7IzUzE4ZxdEEe
TuesWpZUp77TQOu8h1wVRmOIfu6b3grbUik7Jet1cISBZSvWCaNPe8MwiT9audC+NXW/vJ/XbbDdjEf3SE2Hr+4nKfDziAKGsyuUqz5DVvxJSKoT6O5xjvfYMugy0nzD
BmRQ231rCqfSId6H9SiTZ+Tm6hNXIK7qnKN6kLDvRD+eE+puhSfZIpM/lJefljVq0ZaNzMpFGHxUbdSpKjgBCuaqK+V+cA2JiLsaa6Nnz20RtZOzBbT77uFcEwv0sDtx
s2ostqXjm5xsJC64/c2F3cvpZf51B46sqpaaglwhMWZw1JQC88nKjBG+0T3JYNWPYpw1xRdrqb6I68WnXEXwBF0aC1ymFWWLcUN0Vs61unBj+JX7iy9zJTrAORh5YcVE
h9gCtLB8wLrul09qzXZT0vJDtuiTjcHNxPkE2bEma+zihCLa6graAOWNbEffSrIwbJtrqOiqpQ/79gBy/osfUxaP2pWopgvtbi+szSlY1t7hF53yM43iAa6aGe/4BotZ
InCJMLrFHMEsLA34LQ+BQ/Jj/1/4Tjn+Txr/VwilacblimD6WU6Rx1WzVRifwWc8lBwn3BWfE7l7oqqPzXoOaskefiJ4rz0+1xlq+1887XpwLq7YWyn1BI/vmp/tNX28
k2zKEjREFKnVvxsKLmbOz+3Y1/io2YGpgNnS4+7srnPRSUdG+FSyt0SMUeo7fqXKo2qEytXsjrqFF1gCsPzv5m2mzOqryblg6JDHmh69cjO9nl/gPW25ON+N38P9VJAH
mBOWgFVb/zKW/IeyQobb1VrGrklMKvHCF5Kv34J8MwEc09W4Crb5tpWj+ECuFKGrF4KEkQuFOzPBMx8vZ3dn0YfoETIDLF9uh2UKKyrsmsAPfXjL+HpJ6gAj7czs4U+3
irIIz4hpofKvkWXCe+QmH96QkR50Dc34e+5d0X8vURHTvSk87cNa58lBDStsWHl7mCj4VPik+n4yI+Qkt9/L5IZZdzPbKyBztEOL34ezoEMu+ft0c7XjPEspl7/SRVZs
4dt9CC4r3tRfHTFfFzv5/lz7ibl6RKSVg3lN2DGn94SfMMHIMmBKmJHW48iH7j4LG06ePao7OySi+WRpi/X7pxOR1tQXak3lqp3JY2wpAxtVFFkKFDieim1roM/BTgVO
EBrXnx1euiQ6iHPQLHViwPEJ1Hth+qlOGzffbE77dHJLwVQvryaKUYXKto9XbxwsZ8iignrjCzFcBWrpA6oloqOJMBFics+mzUizKOh3TrnaslsDb5nuFcso5xUw0tU+
DF4wtA/VVfshGzek2hzqLxEykrvN63EIB3MwLcY5JQIHYF4/7N7y2A2xaV8OFAfkFsz6xcrrInt5ZAtDm9joaoOBPKQB0KQgE86TXvO0KMa56E3ji3bAeLqhx47RD18R
5xQ2pu3cYLSW4LSW7AeLRaIg0lACDeCeTPXOqpupJvXuVh+LxQnbN8Cw3p0OYV/YGjO7Nobifp3RURp4u/iY9T85oImHpKU9PePVw0ukGwwez8j5yop+miuw5HBco5iP
ywaMmq7uFhsSH1BZA3+j3vL60E/yDfasvCMWvfcsjQSGT7/6rgc0AHrmGZBAtBctYmS5lVCg/ye/zlw1lXn4Tzr/YvZpsXn0e8WdJYM9dcXXjpdyZmMzSKr/LUyk4qJB
4D3P3nwi4sjWC6azIlKedb38XZCBXzTxEzBCaOFlUOWQtWQ+4CFXjapAu4BE3i1y95CGrtENUQq/zg8X8r7YDOQZ4UhBQ8X9lTG897vfNxqZZ3dZdVUNa3ICllKVSC6Q
1EsSDVOjqqiJ9IGXGqc8KsZjNVjd5LP3663ooDuKi8vRczZ26UpOJSVu7TKkUEziRC8+ddX+I3qqUllzJ+z8TCYSLimh/O4F+nDHw2WML9FtpQSCkUkKcmKxQF9jbRtZ
WJRny7n9a14uzVvQEheVn1P0jAeM9IZXCvaFISlqDuKbuSCwP6hYUKvZPDM2uAYw11U7hgGLJrduBnz1cOKsiXXt68Pj5Irku4t9IYgDN6ybswkzjezodUU2FOntDZX8
AvxGVp45f9X3WFliQvPCq1tlmIh5Elj5W2yrJk0j1PwMaHF31vK4lsbiGoc05xuQYVXqovPBWzVooJNF3OrpwBB1Cye1lpS76R5m93aTFEhDAPzLVHaRVhFXND/4NTsR
9ccbeyVAqDsRdftSqz31v1UUWQoUOJ6KbWugz8FOBU5Z/zf+Jm+4Lt1HP/5CU/xInY5EZoABj//gUY8RAQxxnmIkcDWuAKyZLVYh/d2voZPQzAo2GuNH8W4DwuPA/eXo
vgF19ASTksfRw04G3t+tawuDt+vVJF7/DU6F8mPWpxstxOAdXPZbLyBEE+arZtldVOOIB/jq+XV3vFL8h//GBSuH06ZPVHmZFow/V/U+8jLuv06ze1B1d+YWJgHqREG6
4RMAeG4fhaLKpXfEcesV5pn69cOAusEJNw/ajGu0eFZV2v3FQ8oqGulkT3nc50TyvWeFek5F4C0YezU5UgjN+T6lHoAFHDEr0vJCJaJtA0jGATg3CHWj0U9XtrGZ5BnV
a/DQ+AVVqnE8BxYerC3ighvFgdsNyHTQxM+rCoGUMfFnoS2yCyjn8X+tczWVTYApF3WmUlP+cKPfLWwzzG0/I1UUWQoUOJ6KbWugz8FOBU69aDoLTWS65HJ5mk9TZQ9F
FLQ7JVmmzhNnijsCP1Mea8Q+D5NpPVWhdgGZV3+rgW+Nt/g2o/uT3E5pHjY+3o2QPLiqvjJVkgIfmebfypjN9in+ao8i2U8Xj8/okuXitqHTK4nIvcAAjIUrW3rSMICE
kLVkPuAhV42qQLuARN4tcrfVF0cRbN+8On1yKZzVf6hG20GcpQlYMp2xJEVWBnqUB75tkjfTBQb4+Eq5ZO2bVE2QEHQhmJuZbEzAXV41dvIWlAngL+o7xqs4f9NPyuda
WZpvImNsuOBEsoMTW8NeZ0tUvd2pl4QQD3dMXJPpe2MOcAe60zkukQlEWGtGoZDYHFfhEa8nsZJ/jXyFkyBRxJ8+ab4+sBKwxfe5y73f4X0qkd1WRWM6R71N3s8D3O5k
3T7TabaKZc0ivjdk7ygcmLS8o5i5pu6p6nRlKo8g09Ryz6EI6rtdpziTUv/uST/FQUKpn8OdPs5lklzIDDaJLuYHakC6K0laCfT7FN+qQnvlHABZx/SooGxeQ/fS50XR
j1La2rNy0BElz9dTwufSoX/ET9bx/Eqgc6xla146AFswC3q/YNxF+eMx4ZYT3YTfQTSleA2SmbrlZtKT7L9T+nMIpdihfdIRCui/vXdYLYCScYQ3ULHWeSnCSCc5bQXH
SqgGj2JGMMKqTg9ULUFiXP5Sko0szAxVD87eus+20v5USdAh31+Fjm1g4Q2IhgQxA9E6sOqameVxwJrCgy6MlcomKroata6pXbSDY3GjTRCDgTykAdCkIBPOk17ztCjG
RFvVK0T3Xboj8GJ6xGWOGz29jZIhuzkVF7A595u2G8+vLoRnKQTcpaMMjTOytu5wKvnxjQIWJ7625vFEr6ePpRs+B0PbG/u73L7quGn0XwjzWlDPY2AOy+fWji8Y7AGz
4pg7lMsb9UVn+H/fepV4+UxvZQBNw3rjiQHAJHeo2YFHLbqRE8UoBt3qcaLAK/DaMqLRDyCOcRNojiz7w0DhP8Fic7EE49KFgF/LnQu5u/iHpEWVRASW08NmkmicOeKS
ipzXM9SfqARHzAo4niufwvVQRF4wU1TMUOfmiJc4iLjW38U+BIvxaatvbphJVQRBIwxHE34BnE7BeUAEbcE4MZ8+ab4+sBKwxfe5y73f4X1ki9fahJulYRWW33HV8VKo
HG46MlK7DGT1ESxJhgrd4LrbZ8IFLjGnjCFDmXFh17/b2ux1qj4k+SdXEzdqkCzLbVxkRYI+FBS7uTD19vWT6mPKGwSrgg/SdjB0ibVvnZIUxHhNJl5wT/ev36dFR9o2
+/sE3ECpcjAEAJxW3pzulBs+B0PbG/u73L7quGn0XwjzWlDPY2AOy+fWji8Y7AGz4pg7lMsb9UVn+H/fepV4+UxvZQBNw3rjiQHAJHeo2YFHLbqRE8UoBt3qcaLAK/Da
MqLRDyCOcRNojiz7w0DhP8Fic7EE49KFgF/LnQu5u/ieP5OU0dOC99+l6stVkZqBRIW5IZvtX1+jcXdhWMRdpfVQRF4wU1TMUOfmiJc4iLjBxMc0OKh/vmlevZ7gvRZC
IwxHE34BnE7BeUAEbcE4MZ8+ab4+sBKwxfe5y73f4X1ki9fahJulYRWW33HV8VKoHG46MlK7DGT1ESxJhgrd4LrbZ8IFLjGnjCFDmXFh17/b2ux1qj4k+SdXEzdqkCzL
zCKgtsIQ7Bz2ba29khWMYmPKGwSrgg/SdjB0ibVvnZJiXKmA6002azgyWU0yrZ3dUEx/fyrA3ax3/X4d3ofY6Bs+B0PbG/u73L7quGn0XwjzWlDPY2AOy+fWji8Y7AGz
4pg7lMsb9UVn+H/fepV4+UxvZQBNw3rjiQHAJHeo2YFHLbqRE8UoBt3qcaLAK/DaMqLRDyCOcRNojiz7w0DhPxKxDrXkpg4lWA9bLqZ4ollAHz4prRPEEHvEjQObA61g
l+2IgWMXWjDLCnxkQTxg81XX3RO5OSEFJbUQydfw7OTGOrpPIKvsUvJ0YEGFA6QSDi1JAM2zXsgRhSmvEwzn//Bpb8TBsR7oi8L/5PHraH5U44gH+Or5dXe8UvyH/8YF
BqfOTH7AKNbcIgNmrRDpdR7PyPnKin6aK7DkcFyjmI8HVyQNPdEOQd609HdHBYsUCkyVaFp3qAUS7Vsgp2W5t8J17tjfQW1pglH5d63Y/eTEcsjY0wNcP3xeJUXHskEb
3+D48ZhENEx/pPhZDc+yGmCh24FwV9jHRPvprq5CbOdEW9UrRPdduiPwYnrEZY4biFfHbrw/SU/SMB9YDnfFGa6xpf/3MojVHyamsn4dVDlpTI3dyZCzD6m4KHqZ3sfp
NfSnutZKxB6Zb8m4UraWeiLekvvtAkGdIqA9695Egd6urcoNtfRk8oMrQcpSqtl0rsmt9rODcl9PswsmHX0AfuaT7sj+FahC7jeqo6vjk2BRSsjkC+dwtA4xTAEKLZLx
zl1OWbrrM4pOrI+ceug5CDr/YvZpsXn0e8WdJYM9dcVsQlJ3vb03JENd3TMesfswXpS4tDj5xHnJiwgfhACThLaaD7vA9CbRSajERc1UKlMD0Tqw6pqZ5XHAmsKDLoyV
yiYquhq1rqldtINjcaNNEHDfCiNPfY31QYn5KYMI/lhoDsPZriU7R2xjHopa3tvOKpHdVkVjOke9Td7PA9zuZJu5ILA/qFhQq9k8Mza4BjDcoqmnzZ85fqAu8KgURMyp
0c45o1yGTR3dVi0CXNvU+069oxNTVZ4Tpdv9Qv+HTDb4HZWgcjfB156Xv80cdCz3P8xJqzvHExG0AlUqTpz5rx9grJLU+mRVeT4nk/1CIdpmPyGu5EBaYVPgaXsrgjm+
qIAd5fJ2KBBfE8sHRI140j29jZIhuzkVF7A595u2G8+fLb9hNqee2wjSTPYA+sh3B2B4drgDVSYyGdbjgNxd1P5Sko0szAxVD87eus+20v7fp0LCP3wFthAjZ2fD7K8V
nnpyisoa2kLR2fM8aBtdVKYbJ+gD/28GsCwE5g11rds1oiuPkSeA3uFtM1lUjGBNVm7/8N17kBHpu57n4VzH15cduCYYlhAqBLWSWcdcf2cBvIg8bTSb/SKrXA44fJC/
W5OcSXO3LmaRYZib+bhhxertqde68HMPmCNRHEsnB035FMSBhG6SvEpVKV97cIPhh6RFlUQEltPDZpJonDnikiaWmtJQMgp/FiyXruNpyXFnJT1Plri0hSLg+7mh3YsQ
+sTrg3KP1Ze6RtzHUOBQ9qrkz6qMoaLNoGI5gFyohZk6txujopMvF11FAxO/slzYGgAG/jle7y127hJy/g3g0t0+02m2imXNIr43ZO8oHJgYSFk1E54Ge3VcxwxgzV5N
PN7x9+3L524593+T/BO3yAanzkx+wCjW3CIDZq0Q6XUez8j5yop+miuw5HBco5iPv/sz5rM5+aamfo2gNtU8Z3+fOcWUzX8dkUHamAo8lMO2mg+7wPQm0UmoxEXNVCpT
A9E6sOqameVxwJrCgy6MlcomKroata6pXbSDY3GjTRBw3wojT32N9UGJ+SmDCP5YaA7D2a4lO0dsYx6KWt7bzh4w0czczKOPtN62vNTd296dggbWsUXwRkekNk7tKPA2
stdhMqGBkxroWBplnNnsm16GZHDitVr1gzh4YHV5BqHFNfbONGDuSM1rFVeWrBB/MDovZL0otu/F+oNfc9nacdcTtO13yJrER7eK+dj1KQH00ipo+u+cE7A1burZjyB9
FpQJ4C/qO8arOH/TT8rnWrmCRcO5uQkejKcd/4K5ojiCwydyzrpCgHXHfo+AUiKaXUZK6UwTlebo3nBoUT2yF3w0FXqAAkEB67CQ+29lvMky5RYuPDfMVH88plsD08Q/
0kOqG7+zDMtJ/0BvjaUJAh+o16V5Z5JWVN03qdxZXV7+UpKNLMwMVQ/O3rrPttL+36dCwj98BbYQI2dnw+yvFZ56corKGtpC0dnzPGgbXVSmGyfoA/9vBrAsBOYNda3b
NaIrj5EngN7hbTNZVIxgTfAVPQToYsBGbpoRoAsiIMvdPtNptoplzSK+N2TvKByYfYsBdnGzazm9gDDLGDyqocPhEaqIWWLgIKy6+B30b854eoAamCAlQjMyLVQEbF4K
3I9OdBvobSOOWdXwUz3FcRbKxu7J7q9iXbe7t3Ntw/0meaMeS+Q5Bm2xJjSv4FU5BnY18wRjVDHzr1aWthDoWIZ2C+yKDlKz/RTXKLW6Fu8u+ft0c7XjPEspl7/SRVZs
3YdtLSeJw1FjK0/ETxZbE2gOw9muJTtHbGMeilre286fMMHIMmBKmJHW48iH7j4LuRFQ54hdOaPxU9WMIWpn9vaNo0J5QOvPxmZTDX+Q+ZIbPgdD2xv7u9y+6rhp9F8I
81pQz2NgDsvn1o4vGOwBs+KYO5TLG/VFZ/h/33qVePlMb2UATcN644kBwCR3qNmBRy26kRPFKAbd6nGiwCvw2ikjk/2/qOHOXWQ8WmPVaRgvOGS6c122JdEulT7vVweE
XRp3n1cusUx0apIlvlw1jkBdtpdVibgFbYEV0QVMKYocbjoyUrsMZPURLEmGCt3g/AnZhPhIvxY+evH1Ekx6e0hcWwQhiaVddmc5g6xkT4lRjJWuQJt2VSgZQ4Z4Z4NZ
KXO8BlKKY1mIlX2IZb0IqgkopSrobSBE2+NBEVwsovWVP+Jy41Mm3pxDRtHar/pn1QJ4Ip2T6byJ6K1e6weAlF5CIkQZP9+OimtPb87uvhq9pN4pLntIGj0q3ISbGi1m
8HN1Nx5fX3nW1/qr8jU0O0yqnx74jfmHdP8n0R8QS6icdiNrdA67qN0liysPg6Go1qB5mHuf0bn95AvS2yFU7j8DyETtD1g1+3Dg93IXzLaxzl06CB/QsFnZYGHbQBlY
zfSYTC5xthoCPkydLA7zu9XZ0ckAgyPcsUwO401EbM+25oD1Y1V7wtMwGUeaQsNffKX0qgKzOU2CZC0vogm6xFEfn9a4omsZTBnmgibvfuFn+4F2A0jce7KrgjtIfMCH
w3nsGJqVnIgY4zY2wHUXFLQaVxqsvrB8CypWZawnYEztIkS+JPsXLrXq2ebSHThG7x4dwZjRR1+CrGKnDx4a3255Xcs68FWbte2skq41w5iO3a6KkF1DPPLWb0vUBhjD
fVW+loNk0RI24r4apmoWdntY9+hHi5avNUV03ZSSzQSgwJoJEqGByzVJx5yqHK132d5lj4Nu8KtJ30avSUONKzfEE8lWwdDTXHsmWS2pmIeVugnZf9BZSvjjpcr/1YCv
RXTc/qHI4jBRMOj49YLx9rVDxmP+R4ZpDOQPHyYvFHvTR4VCDExa786K6gfccMq2MQvx8lbibNeYz3yy1XAaQoI6MCMe3GBD/ID7g/wQNAiz4MKbIEJIxRMhEND1mXqb
tk1VQjbau18cybdzE232c1RCzKfEFLJfYywJMP2ocopTn7x8n8PRgHp8lSh010Yl82FXGbXEw4jatXJmnJfvEH5U5mjFoHZIAOcio8rNKUQ2ln5cu/4nHVKdD6P4puaU
LMFzCO39jvX4q0U4rF5pqYNNvUYcHfvKV/fKCszOhMQA777TbXbmC1VD8g8JXYqJRzs7ZlKre+2PL0UM9w6kegg6CqpCc47huGbu36wXFyLbuSJFwgs6uLxAL04INkPj
uM690pQunEZpGLNopI3fuxWSAynpHCOrCJMDeiD4LENiGtPNZ5vmCO43LwbMtUcNl8PvTxtL8LwXI9iphZKmhWOu18JaaaFR4oh5DpuJxtZVaIESn1QRX03fwk4btO1u
PMDR9+3dEoW1jwYmAKpgMyMrYl89mSPsbEo4oL+exxYqYa6e4F98wJ8xoAo1e1/5lEmoPEDsXWUXPpsowUnn9Hx8enMUPy8slrJzLzMbHn7kAU7Gnq21yHBs8xzYceYw
sqkJiR72GMe8+mKkAyVgfAY5BrBhB1tzt60e6SFfxRWJA3DwYSpA2Adcnq1L/+9/rLmu7RZxzTHJwRXiYe3RnVGJuk3/q9HFJS4CYWCBplK1c5YoTO1AiNL1tfiZp/sZ
ybrKYgFzfWxaxF9xWlmGdWY3hhUdlveVC13guXiZOzZBCobs+zCLOxQ7gFf7CU71hdxUAssYHKd42U6nfdoD9P4b41EIVSF6WHHBnIv/SHoJ4ACgSkitPyPpyi1pHi6k
dKFi2hpq+RsED4dZORM2DdqLCAYHiDEXjSJQxEvDDOdf08j6/6/4pZuL0P2OoxSt8aKBIokaKbrxqvLcSWECTw8xf8fSlhX1p1AKRoXAWgJlS/h+lm33mqNY4G2bcPRy
WyD/ExPKP+F4HCCIBNYx3/3QjNZPf7PLZ8Fauc53HHDGw+H1rLGvQcsNFQMrEJvopP07eekv6CyP+veSElvPoO1KBRoYy5Y8rsTzxulTOh3ebWGXuWdJsI+8FhlQfq7Q
6n2ZdaQkO0AzKiatGlqvYufKB1rSLhDK12hWdX0aW0f/BktMGvJkrOVODlt+x2//Vuk55eNyfov6RWAM6jZQ8B9UcxK+yunDqBpdAvZ0i3EAO3VuzL40DABu1RF9fHyr
RvFhMSFvkQm4BQ5nyOznXR1hii34N/r9wFSkcLzvQ84LmKGG9DmLNNO+q0p0YTEyr4U6NnGIOvsGsXLIOTxxf/A1ZXEkt/4d6NIMKtwxXNMP/KCCVyqCKulD2XHVgarD
iG9t/Kj33sCUV46LvPQcm7FR5IqN8EpGBvYzBhJ0CGw++KmW5t9KigDV/zwTwiMZaXlkyF3TYt84d8cbwNsWte0o251nZnN8FyPSD8/pScN+jhk5mCkGMNf61zE9Yp9H
MoniPAbD5wCaBJwKxESG21LFDHPM9zvWILPdElF16IKtkJSkiMbjfG5sCjDOtiSwBtwsI4qbZa08t2l5x+jzdM3j/TpMLIBrJOgTl/IeZ89jInffT57SrpYFVYnmsEfw
jq1gRTgIiKNkfkXMW8tBMbLp2GIYSVr9TFK1BExXTAbVtrGloGD6s1tlG7/XBANPfxa1rjDlcC83Jt8t1R6qrpvP3CC1209ORlaqsEKcWLPuchyCOUOHHTlI3+v3Vmld
0AzP+OTYQVWD/ra6nbkZt0VS/CD0ROnV/609ag1qYH1pFDNCcd2pTSYYRqoC/rG2ZO6vgK8ZE+r2NOKlRtrfH/TeEjlsqv+F3zitm9B/dWA2JIBZTUok8vwxEJBInzlT
TTA7dkIO5RdV2FI5TVPguQfbcrNcIUwx0ygqHpmRMBUdg64NVYwg1Xajd8fqSRyYg7nV9E9H3t+bQoiRzeAd8UzgFfMddCApjH4zbJ/kfcWsKtyhoWqnx7GxjNqR0aI7
6mk+Vms3WOf8aHvfdneWSHAunZxsyTK6VTocUU4lEyZP4X8gulFCsftFR8FpPUbMgOAwGp3lk43e1S/6030QAuLL0RkrOXWu3QhG5kSS9YxjFSBNl5qFo4ltryt5MLxR
U2eg7VEhRJXTvkNe/trjNlmTdvrf5p2BWYpjFI8Gnx3wX6hPHGSFd7X9uQpmNZ0yOllN51uTtl1VEkG9U8iPlHQUBkECbKTGd7SYeLHit/lNsA0/7bnrcAPDtlYWYCMc
x7JSOYsNS1T4e3tuvv+DReGAdz/tURlxV1yeem+E3RyGoZFUTmqCAXv8zjvIAs5sBJVQrjYOZCIX+7O0lkXZTLflTO1UCziOQk5orjrK1NxVaIESn1QRX03fwk4btO1u
WSm1Nj6w7HlNLaMVNh6KkVRIDxBkNLStUVfbNOZOaRKp28vDqsSpHuE722VofHQxtyWq0fznl9ugdhagHX9cfCniJNUDS4ny9F7ttBuxeI+vOjr37agMDkbC/shKSP99
x4GE31VIfLr3mRHjCevBr2+CCtECbE/N5++8ZSdy9NDuR6334n7vBc+uvtP5jh51PVJLu99Vqc62czoMgLEyUfSSR1Iz4NIxuQfsXXsI8Kad4oCqYlY4e7I/+P2NIPsS
DzF/x9KWFfWnUApGhcBaAmVL+H6Wbfeao1jgbZtw9HIDb/NJnbkC1EjV/1o7zDYE6U+/eeFV+WTK+WfwYJYxmh09TijzXxIj4djf5AdjUSFLR8fUPch2O6a2gWQkaRv1
6VsHSHWETu2VpzIqQbMs1S1DwsEoM/V5E5Ms9Xksf8luSs5tK+Ze2G5o5zNBKG/ljU0Vbj3sva4gHPMQC3Bg6qrqKg/0Jilf76cO6b0MC/RsiPXoNCjJCbTi5IFDCNdO
od3kTT8IKKJsJbQ+jJ9v/6VO25OYKG5WyYiJ89U3wxjrCiKBrUJJ4YZVNX9KwYGJ8igpivyDPevkmMTCiTCWpi/0ggST5KZ34yZzTz1CQ0HKQ8R159LH9eyn66GgsQ4O
ibXzAZ3+ql7r4wOAP8m8gu30yCMGr7IIPNSEpfxugfMvioZPOuM3pZSqCRNk54CvEqsovEh8khJDYhHO+Gp9Ry04E7ot/qpd8ueVUTNWmUf8a9fXB947D2ZQsCajUZhb
HnQzUXjHxQPFyY+x2snAn3VlvxNeJrykF3Hp7mL58WUABXww9ZJr6Vs/M5hRLRQVX4H9nUwKpqyDVO1KNExDLGqNNX2XTeJ15THXL5qEBjdu/GdIcRccjFArKA+gecO6
cHKLqXUHF+sMbQDSBjQ+DYc0SodyWlrFpO0gVhh8js8nFQGFPkCsDG9b1ESzO4o4x02SizZMK/oNC3AvXvFZ0XdLat/wPAmsbcySJ1YiXZdzmSgfIXHnvZr++OloUViY
zf38dwGAJxwV3X9r2PiaiNvg2zoB3OKLeuJK/EgJ9M0YNNxXVnldZsARgdkP0HuvYudOIoQDJVxYb+BRDJXKtApPY3XLHQIuh8xBvTKRPRD8LXw7qC8dcrmGGbbK3QdY
X1nT/xS9Xc9oPQLEdJRsJVS3cVTj7wf6fyVP6UXSWDaV1kP4qMNg54udS+qo74Pat52oxkmGLfM/tkXEdX9+NeFIWe2ZG4/BpuO1JmCt2WNqTPNu5AyuTL/U92GbbIbS
Te2OJTDKwVtGR5gobKpBq2p8Q/ap4fqLE2zE5FCF1r/+gT7GKMRDkoW6V57PsX1abRVIywmaeJlcENTC/WZtE57CQv5DBGcEK4D1JEkQwyr2gTqTwOApwJW6Alotxcu6
ez/CS1bEzQdzBZGyPhkSTlmtz7BoufipRQphLC8cPd7l4PRxYLtdCtlEIpRTYz+2GMX3PJhFxPfBjk725O4MnRPx+eoydDKhLb8sszOpoKcNbFUGVeY8noxj98G8UVOG
kSUwqZkGzCPAhQ+Lacz31hMPnod0EI/+O2gnALWVQZYr+4t5WRDicl6gBvC8hN1+JKoroVgMeSdDr8ysymPSCvJJywM3WoP+4w7MDfF2ZDGMoZTRpEgQM2DK93i0OKUy
0/Z3GMEqCEY9SC9KBRANfyBDzw5VguoqRTliybLUOQTkZkyhtDT4vqYNzIUT9Vk5IQoDFxWORtOtnascjIShYym9qqmXIEhREUaCRaDurUHQBiSqBtYo9ZEfFJWG0avD
HNBG8Cbb7QmQZqojQCtLXSlBACDIj8tWHBYvY5YI/78F10/eoTtCFfNfZR493IzVG1ubSv0y4ROyfvazLLqfsWAwQrqR7uQwXSrHzxgW0cZUTcPuC41qcEOW/c8d8W0I
PO1KgIETx4aeIsY42a1bKVfhgLWOWijvj2kfJEagqtXm4IQ2qwyyMXppgk+4UaVT4t9p8q7FYe4++FEy9nUKziVLn7c4i5G2xxviyFUDdWWnq6/keYslPW+b2bGGjMAc
z5nFCYUq+QWcn9I92n0OzaXZCbdL+AMnqSEq/TwKkfSkm+Epzt0l8fxmrn6JJKYta+edWHIV4kBPs7Ug5KXHd6hw8SfAeNT72ds/hzNGWp3GnaS9v/WuKDvatrrqCVrJ
fAOkZiQUam96YD0T/Y9aNgHZ+Wt9882KA5zT+LFFQLM0sKO70qUNbyv90Ou757V6IgtXIMJUMBmgwY7WFp+rfg7+POlfqX19ynmVaIMxrivwod+VpPHZg1FWZ+UP11ql
nncLRYUETMfu8zaqlkKBDW2C91JfteIUPHss4VVI3srNobRJeRzXTlyS3RXYIYixkl0vRQM0YAMtS4CzVIgQv4EjqmK7AAwL7v/hjPcAyT0r4EqB1cEr0EmH4y9Wa+G7
qmutStkTknzy8Fy4uiuJ8Oq8GzPsrak1FQeggen7QoWWdKiN0GYB0fk/x8/FVnhm9/oa03cIdvFX/s3qual480upP4d4KZpDJfaJn0Wno9YhQ66SfrqyMfmhoo2r7/pd
7li8OZmDjUakXulyrge0X46bbyq8ZzUKTBkpwsmUadQz2NKb1amZzBOdjFfNCmA5dcsF1qm5VHw5rnrzUuijruGAdz/tURlxV1yeem+E3RwaN6U5itYSVQmpx/80C4w7
Lfb/2oK0RRUrF4VH/BBAXa/up5ttEroD+mf/hhOL/vzMNijukMB4MSgvj7crxp1eiXsxjmEVW+IEsTtcnY5MWwzW16DM5p8+OXYM2T6b2L9G5JWtCRRUZGXJRzwfVgWG
dXB16jO3CSi7k8b8Idnzmdjx3U6X2EfPBGNaH+scs5Sl6LR8EaUpLugqRDcOOGsBShk0BOrqXMgMySJMFSSOttjx3U6X2EfPBGNaH+scs5TOpqhFbeJLwy35d8pK1qKC
XX77wgD+y0eJ90Ke6YxDiNjx3U6X2EfPBGNaH+scs5Tm+nScCZxNp3FUGgC6AJMoMVRLBGYL0ope/4ofrNI9k9jx3U6X2EfPBGNaH+scs5RZwXSkYADNBc0rvV0mb0+O
GI9imePOy9Qomsn+vPVvyzo2s7lmrqreOmwElkINI22gFYjD7IHDy9ZVoAd81lankBkj2ZZHFsQtFjTs/OTOEjo2s7lmrqreOmwElkINI22+gHtokS/BSfI/02qZnXNw
gRYWEOjiMzPHp1Ayqc9J63ujbZdki42miFK0K15sBvJRtM/jGSMoG2a4Z6MofSk4ZgcLIU0Ui4AhqfEmmeW20ST+eRAQfkaS53JQ3Yz7him5eMA0EUF+YacfiTALmmkS
ZF2Md6q8C+J1zTvy6Rf6jgOWNbsAQWhtTQcD7hH/dMxq2zROdew4M2wzIwQRRSgX7KeWX754RAaL+ScYYUqLBdCpN++KhExuZ4IIfneWGigM16byx75Svoqn1vEE3yA6
ATt6SAV5Ruh8F2qJ8Y/DEKg3qljP2NcLN8Ugzv1kTOzJMeMuTGvG5/nTabeCV6S6tJzdliK1/Ql83TYNAcSYFOUailte0ZxGgvYzNRUCuIoWaXDGt70XzaFjjGR3Rvf6
PCorEvOiHsiJKXOhW8oN6O3zmdMohxDmBpN//BVHjtpU2xtJ5l0TAm0ZK9km1YTVgxj1FpHBfvQgHSlVkyz5od72BixFkKt+HXtlO+CWLi/ql+NlNQHGVupYJjTMbWuv
8S0HbkRMmFAnm2RxacU7O1lyYP/h5KGdRdmJUwrj0+233qcF+p3wV8oBMxZRAZ1F91/IRH3qCUfOSCDlzI5ubNO+oeBXIVxF1UfZJlNTcNbzcQClMob+AEeD3P7jqtwi
6XrPoWbLNVvuLgP3n+/PcvWoCMujrv+zdmB5yDv5IVTRYVKung+ErL7yFdgS9Rk/a6o6SlftqEjsHJzDqgfoRqCyYfTAVjjOSkx2k8EBOF+k7jBayCXV+KqVgzC0+oa4
J+cvmWkLg4ixMlbYf/OTfY0c5Mary6N5FJoKOku67yNcorTU8ufmVrr6BSc3byF0qxNeayvwLotUXrsgpkSRETV68yJqrD6cZ/nSv4yth4GYVD+i7AshWBcQfS4GFBZe
VK++BFzsNL0OkjuIQ0FRtUq3pbMeLVfdmRJ6KXtf/urrFn3dndKYRNkt6gLBNdrdAK9Rf0qWCAL1ZDe3jPV02sgf/+U7DvJLws3KX/T/dYaLS3W5bYxrXE/wCEaoQY8J
+5xfhqu/AMy9IVR4z44DF1c3RYOYO7foS8irC4uLWWLB5ojp2PE8wWUwNZrcs0U4oL6mkwfgoSqIC3Jx2MjwOx7KwI9XWyB9ynPd9kyAZLH26n1FtTnxSau46N+UKhCo
wKOscTD1T1FjlG6kb+hFQcqGHaCnUQ1BNJSevaFL8dzEeS5Zj/8usOfFGESJzl3hW1pDRIY/TKsnTwECvsGBlO/dBqfb8TvF8S9G+/QZItEryaIejMiHbfO3agetscAR
6KhUQ6681xje4/4xQn8viHyCjT4LL7M0lH3AxNO1meM802M4j18ypDwPBZLnE2TSTbt7fPlJhX6rJOyo5lFFVt7Sp/LnDZ+sxA6IPdvMf5pOHnBpW3pjD/7TLEBpHdu8
c2vImaZRXip8Nk4LGNGDbNamei97za+ztn+Yq4x39sDsklqJL3k/do2DuRQ/ceKgmpDu3zCEdlY44Xew2vNxWR8CzjIHcM523egwZ1nJSIl14XqOaPM4Hr7DTvUmp/gy
/JIYbD3a+1rHW9c57HG76oUW8d6AttGis/GYrx2Ktomqz9k+3lqyK4bwONWVKt7G98DQWYbKQk28nnBuKtcRL5+TP7/VIn5rUALcOR9fS3ATI+MzXrEji7rJ0iW17iew
UtubGxRmjS0I3Swpemi/q4GTd8Pep7H2w57Mcc2ukwD52Ox5CDg5PuwptFerSSiqoxK9JUvsxg+iLMySIgiLH0nDNf3ntgJZeXEiF7ZuwWXYKwUbfoViCLQRHc6DQjjA
k/gDqnM3SlmQk4CTCktsQNCT+dPdwjpZq1iyCHN6ANDv/YhtBhgvF84eaYDInBXPpM6pUM+1qe1WH9xo2gWrDE8n3I5Awv2Q29EUuyqChJAzVr05/u9SZMnSCug1DWrE
8kHNnv3fyExdzk2QNF4fMBw60EuFpuMBAUONP9uDFUhTB+CeMbkriyF266WkmwvlVJd6QCjeb1XrOEzsziWLLbWuaRLSXxjuUS/pXVEX0+rhgwbH5G3VjjfwqVsy64Xf
mxBBLG6tUpVeghmnT4+SC4r0zF9UdQ23Scxn7jfmqMR5iqzYNfkWsfsSAlmbTuE/lfz8q3niiMiot5tHqULJxbryOUhchXgt48h5/R4D6UU7EuATmycLCdgqYEbjVquT
4G+fYMi3o+ExxTgZzIRlPJ8ucVGv9PpDcKxlzoAH5v+mqQIe1DHfDck6LNgUCBVihzazGbv66InhbGKZks9YE/0RKNHdTb5mQFvvj42j2Ffmt0TUYkJ+x5rnaD+yCnMA
5ObqE1cgruqco3qQsO9EP/dtJjTzEeRKsW9LPPEaEXs0bKGBTETAmmU2o1yELghCtNNqkOkI3OjoA0KJfScoqetTYvtwW93wlJqBwIDW1QRP61yuDnYX2urvFWb4u4VT
y+ll/nUHjqyqlpqCXCExZnDUlALzycqMEb7RPclg1Y+SmAWBSuqVAxYc7yMfFa5GZORFiDQVAjZQwwWTjE6FZK1WVPtolBOFu4qPRy0+0zksD5OXDjsMmxU4l3FJRlE7
LGOOlYDveSXm4ybdyAyYd4yoFQOM6+iBfeGYRwV4BbTl+m79U47dHIMzHb6fgef1ofstrXX5t2tJlTmirjhnUl8P1BQz9hkA+ym5vQRkRn0ksYP4cmzhGgGcOhaEqfvW
BA/vS/Qskklyn/fqoxjK7crvAElb7OBizPFg3IJE4cgJ8sQExhULfYyWzh3+sNgK5lUBWR37C8RqVGMkK6+WhtYdqzXUr3PX2V4JSiWaOzurzVciQPzTF/0db0RkO75P
0uhNvMSKKyoxENLiCOanBYKEaGR1T87kLMgxwg208rG0rpcT0EgE4HH27kwmkTjdq7kmX3wWXGyf/RbByJhKiOENNSkcsC2hvE2FfiZHf/27c+DfvRWdXuJjX0oCe4L2
YyGBHaEvUygQkT8nj9nwD6yKzby7sPO8ErCASquhVHHGS8md56+DpEytEkrb4KKwsh1IvZUHvA1TP3AkHOg5cU4YtwMMGFuz1fPq3ja2LYf/ZfkAZtNilrzoKhgM/htT
EBkKTWULzbLvojosBCZ/VY2XgXJD8pW7jhGGlc3tSLkbq2vIWw0ADQG+omFUIbx1KTivMXRJD3UwKXUekzFN8esG6AQ66tQiUYWIB3FA1mIGHsW9amPul5wUclFWHQL9
cqMrzA+exZ1bvq6nD0PT0Ua9XneHqsRh99ZgoxSufmntTv4mSLtWsjGIpLeYWtqfDuXh2bRAur1DC8FoOFdYPhKxDrXkpg4lWA9bLqZ4ollAHz4prRPEEHvEjQObA61g
Yuj5UdMU7sfTLiol60hvOkWSubGPZ95kn6wET5CinIPUl3GRI/DDZj52PP8Z1+ZTp28pF4KFuXbBZD/XGWZokquv/ldNm4TyWyXrMlYL1OrTtdMVRt04FiMbIw0W9Q1j
h6RFlUQEltPDZpJonDnikoJM3azAHjX1eTeRFvag7qah90D6JhkeSuDWIst7D2PsaWrP/2HDk6IMnnyLFzHTIXQ2IHksrYsbeh2jG05Rh/gwknYtoH2sF8s4K6iS8rX8
U6GTbLwDTr2rfsKmFwXDoiLekvvtAkGdIqA9695Egd6urcoNtfRk8oMrQcpSqtl0QvToZEJXyJqIL8eQU2z5ApQLSLwWK2r5uGM3WhqyGL58tQUSZnVLwnHf4Dd6nR3a
jIr9CG8FgzpMdX42ZWZEH82X0tguaY/boSqgKU3ysAplH/WS5ZKE4T2pS1W+JxwCmt5H118CAbAMvjGG2coqHz5bqqcA7limUajBmqmsNq4jAsFcW+obUI13yJuGsg15
K4LI6R5sxXnCyunoGLrcJG+PfQ/ZjzYLjtPai0Cqr0nDBcjt5pGcaDHJrEqw8zc0Hj7DScC12kimtwtgi6CGp2K8xYdBYVeDpxin8znvprI+jydDS/ysgEfEazHXtkrJ
MCE/rdp4Su4cgyVVNCvoj/ZvKvT+E2JgGosnennJikeQAxTT19OlR0Sr0+SETEJzhAPuHayXfl7Yzt5Q7q3P8t4FnjpWYjiRlMWeBhtvXKHGOrpPIKvsUvJ0YEGFA6QS
siqAzTu2yuBh4OZ1p+5VNdYSuaTiXnvynh4IeY6NCdhto9fVAKyaI9hwi9Xq93sCFLQ7JVmmzhNnijsCP1Mea4ZgsZN4d0lk6Ea3UyUSaE5u1yKzydmf+ryTRxOMuWcw
7KaDSUpYz+7JwOOX/tmwOpj59/X/GD8ub7DAn9A8RI1o7hKVdp/EAv/4dINZty4Aa0avyX4b1IrbIEkrlT+Zkl9Ipsd0un+KfNfb6WtoPG4WcH+9aQj3WaZtlBE9UjSG
9RJ2HkJQLtJvmFHeA/SVYehKe9ZeRkKIYphbQGe3uncSsQ615KYOJVgPWy6meKJZOFJUtspEn3UTJyEaIHt1NVkwQXGl0s1YXPYVr0ly5WoiWbyvmFqq20KDq2ioKxhL
lRbPlhKzp9wdMJNbugzOjdzs2zSYJDHV6caA0+5MOFO4emgvem4TX2hq83lkmelp0d/28ps4zddQHbYcaXJ531AJ1LpMJSo14wdpnOi0nME+1Nnu15WrWGlS93kCC/V1
S8TZH1VDCED8j3O0uNWOG8cyWRKxERVex43jIQtBqHSvhmZFsIMT4hdwbF530wupdxob7xjyL2s9Sqjt/+q+TBAz3F/MCyRs1XmpPf74aySAiLJMjFOag2SXEvabwhp5
zbSzfRPrbHHcXmc8HwITj4Y355YbIs/eRY4iqqEhlZeW2cXsKEjFHM+BR8Jp0sNqq7kmX3wWXGyf/RbByJhKiHkzacBrtgXYIynU9xmD0cOnJ2Lm+PQr6WwYXSQOv0n5
1cglpqZhkiAV7Wio0BFXzlKBTsH8dZojNBgmZrVLzFl3DLifqFv0WtH34sksfHxFtLyjmLmm7qnqdGUqjyDT1FaDd6N3ppvnAR8bm4LIPri82Qj8MSOwNoPNV7osAqKN
2rCIAzCuqOD/SKYAyoqQofaNo0J5QOvPxmZTDX+Q+ZKcAVNiqbsAb6MpdmhDgtQRL/izYjU/VxIWoDWPIR4JyJm++dkuBmsYSvsr0vWd5Z3GS8md56+DpEytEkrb4KKw
NPGGHKF7d79Nl6HRYogg49hvv1XyMMAcpOU1Q7VImNqKCx/eJbQDBmWp01G9/Zpaypjwcn64mDA91JsNy3+XXy7N9TePHnAsf/q0O/CkO4CigeMA2NLOGuOnWWTHBCTd
AdE9ElkedlELJl/hJoJ/3dN9h5bVeIfg3KUoZWsDJnunjxVv4cbox79XE6NmOZJs5wp8A84WVV4JR02Pxm+5Bf8ei4TTu0ykvWFxhDs0B/ymyMWQIMHgGU/KOcSUn4L9
oMVhSv/krFOKNMe95HIMR+MmdOAI/SaWILMkj4KWURHt8mg4OtaKL0UIlo/M3VcEpXBAZO+ch86LC54ZjtYXQC9ZMBf2M4l0Npr49pW2EyQM2uBtJJmoOieAiwbHI04U
F7t+5e2rmR7Y22iGv6UgJGYGVxMWaB7Prn3F/LOCP1//NfgQH5ZdEk56CHxIFfiblRENzKFwrb5sJsRVptL5F+pPW3CLf4PdEuWEVwKlVnFwcOqhR3Sgqcd316brfj3Z
RX/1Kq7l2sXkU0sQEDbNKcNLQ+02PSbIWVj7xDb3irpoV7oprwBh16p98+h9ie5Hf7jY0dwesfcVOF3crUGjHai7aNzB76UkU92sMq758BeUKAf2U/tuhi8y9jhLEvNH
6AGDOgbaM7ar4A8MVTCJGgBCIhuIOTg4/Q9HOei/7DVFpGGTEJLojYMmGfV+As93Ca5gsal+iniG+rm3CBMucn7b5JrJjf2A88msrNdYjP4EoLSLxT6KOccGUeD6HyLB
D6zah3iA8aKXRuRb8UZ5sdN35IxUB1AiSmi0TbE+FMOfq88pUE4f4FvLMSBlst49Bp270idJKORKVJsi4f2n6pDQYGuPy0rZXf08ZmdIlpd/nmYmfFAxpFsfY565xHoz
HwKs8MefnRyzw1ZIAc6vSg85k11BXyyCT/rSgVQwPqKWjFGhAPslvOKlAgSVSNv/IPsOtGCwpgkYjw6YVR804Ll0fvA7KUwKFhtN3iOH9k/UsDGBu8LWY1Ba/iisubAa
TIUkkTBYiQA+wZUIcgdA+DPVSdy86Bs9KecJtnTqgaMPMX/H0pYV9adQCkaFwFoC8y3vTFJE+kdLuYp3LHNTAeqGNtEg52P1kvPiCASPYKnpKf1wE2kDmK2heTn2gVxf
588thNisxmNKM3bU2QhHSTimj1zOicR7bzzyqRGa0lZ8uKmGmKtmqTHi8aFQkTE4mtmzDQw0Y+sbDWQKUMZm9o4Xtehy7jNFOdSCp6fg/fyF46CaDstcQoxfhvoLdV9Z
m+zuxPzDV7oF2bqWszOiYd7vNSvrggoN3RDa1d2VV5QReVfQnCrD97LiHnwSVDn11jjk9HaXK47UMZLkXBTAXHmPAGY5JaNQa2RrOe+v/7Zm4Dmqajr5D7zYkmXFJPC4
Fx1HvyVJlgCfh3fXZzHW/6e/a3nAbpuxaRc9RdFhwXyBpDAsneFB9/YaL8ubmCZD9Xs6R1dWMDZ7LX9kbT7VUflbeyyJaCJUDPAvB1estF4Xb6bQYvUNPGI/vJQdUUMf
PeTFU/9aph/8Kq8kFnep6Uymy3DECSgAHbu37DUKR0Ogj/rYfDFNFoa0p6UHzHxlc0lkj+IrT4+NKbBTMz2j85uG5T+KR9lG8sbeqjLlBoTQclrlqUxOwVLLbVeXEeVp
swRz5tyEnkH3r/ximTSSMh0gzKGYsGhxx3FQXvgchCBpoSLC+FXosfZ7Bs62PGg/2OKCapty+qOdeKZ9mRs2c8voQ/F4A5FqhlayroWwBy9VUSP5nGuXGfFyD4+MiAQ6
UqDuj21NnIThVzCx+OGpWPneycvEWBwvDxd8dwtdO0qTV6bnXinq3KDSuiJj5gd/7Ii2eeZQnC3bAKORK8NkVHvknQRwt/vytjuMNvOHdhH5MV4dSPFPUH9OpNltxIpF
1NW/QDSAMhdMm8DtiAQbBB0gzKGYsGhxx3FQXvgchCAJKXjwr92ZaCUBd4W7lpA4wxIQPrAJm4ZFj0Ezawf4JdoIoDFDsxlVel5SUSgfT4K7qgS/x14BJe9rEjbaC2KN
4AR1req2cOuYU2+ZxWhiJs2K5aSgQ95V+5jPyG+sMoLAsc00IyPGw40Y+YsxFytOfCWBrFPhffV9KgiwyycFy6xD4MGWUSRnk4DsYw0yX8ykm+Epzt0l8fxmrn6JJKYt
haY7uTW1tgO3iwKj6ocUGOKYA+PRcRraLYoTRsZ6qBArRjlTKrUc0VdYNKM84kNnBaX/cbXRjpyEzsY2u27/K+WAKDT+yl9k9kDigB4aZrdIqJwh7G6r3ajxyaD2/xJK
bntk2DgZ8B183k1iuwMGYZ4LcgJpHJyhH2aPRxb+jZpS+tQTKL7WHNFaY5DaiBAxU4N/H+IMlAzO2YeNT+Ijso2N0AAP+FQe0MjpyJPVZx2km+Epzt0l8fxmrn6JJKYt
OADCNLzPii0Z0Uod0aTB7ZbIZP1rplNzT5o771D/9Y/bpJPBL/uT3ysYcLK9YdyNsjq9kydmBHVzRaU0yD0HZx5Fn0oBJVEdL0/Y2LJxsIaQ0GBrj8tK2V39PGZnSJaX
f55mJnxQMaRbH2OeucR6Mx8CrPDHn50cs8NWSAHOr0oPOZNdQV8sgk/60oFUMD6iqenRUXF4gkmDF17zPAN3uXwOQDLsADeFtkoy3oLru1eHFenckEFSxo8/a2ryUiE9
9K8YMQQaYOl6jo9Vq/opUSrL6H9lI7onL8hddEy/aRK20xjwSXJIOwjnz8tkytL6ObKuCtA2n6+w+cgRn20Hd9S5nLb7McaJLAr2fgIQMo1JR9QZ1YSZl8M1Sok5ODOx
ohrE8BesKUkE5/UD9F0cYf7cYBMuzqh5X4/+salPQD6V6e1ltf9NHCme6qhVyQjdF8R2lTXJI1+JqIaVPzfdHyTx7sF97miYR0CT8+DyySg2/qtd3T6HpF3a7ttgALzx
4q1KOb52YBnHD4GHbXRAwuWAZCmxqmnUOEi2bkr5HOk2O77IWHStJN5MY4zPPB6CrvPH8GF9iHDBosSEdDPCt3KTzpsSApq1unXzxDwFDioswNoXVTklM3X8ORpg98bV
QVG2H9p8j0wWerwuCQ0dEB5eKhIIJye1pY7i900RTT5kLOyDATnDEClVRfCDuerdoxkPuY3/3DnD0slu6w4wOLHE3UAwK8F77k+q2THfSEeq5/Eal8wVII+M962/zEGR
zmhHYjYrWLLO5EHpZPREXog9nbPKv0m/MpwmfPCRLqztwQd/NOT8ZpB30FUkF/GAqdl7A7qSXv766l/xUz0+31NsVq7aoK3QIKMkhoboRZ1CN1gK4Wf3iVtu6MP0o8//
EaHvX8emxS3874HVBu0fj6PQwx7Cu8CcLEhkLVF8pv8g6AFurRbrbCrWvGuwzZDGri3HZJrNN+ZZ5ZO38H8f8V8CrHJm3zsWQDlsw2qYC1/XUAcpqfF9nl5yTVAKKRFF
0hYyLFSgxHK1h/fOlb7E6kJo2JOQdDrILIzn7lD4n82irR+OkhHmXsbWr1V2wScLMRGQzkqw6dC0YB9ZAEw0KYBHVi5P/vHBp1ZHK9mWf1E7wBZME0pZl+cFWAQhi10J
xJIGQlTD/zrtxY3bicvJTOqZBlx2PTDllPIiy7hbzUJQTlj47/ixyvsNk2KlE7VLyK/cYIl5/pwyq6n8JZ4OSPRBSqhHnvCcbk14QsKMVtt3tvG+AcX01uwX7xGMynkB
unku6PVEfHpL7+pG32sc2FrOzliAno71PS2OMmTHTPe8zrlwJp6CkVJbsm5LeIRCYJdLvy5rl2TA0trhq835ihl7TckQmkEA6Bkhhpc0vzrhkBCbaEyZzlYRnvexOqw0
o+56/JQopR0/nBU1gTKDIuovCD0+Nyxx29TdFKGEwslTyL/SzGuU35oSETQH/4768C6X1Q5eS7kawHHKhgwvbionxRBi2jg5GKhCxLU8Kc1KXLY9T5QDjG9da2/+7NR3
Y2fDsIgvodl+2Cn8kzyM5H/Oky/IT3XjhMA4mWWAOcpQ9X89CSKANzbtxKy27OOHl49ZqlAZSV/GKIwZOViZMC9kTnh1eeCmefMceSqcpco4xQI+eDvfCLVZAuThWeZy
qitGsCUdOvahkHpxeQ3srqH0SOVXHPp5qDpKzAcBTryFhP2Y2E6NL4FyXxql5vo9cPW+n3OauazL+HEamFHbSgLIjSYTHMg3bv9+Ey4jXRVyhji30BzVCV3HlPeiHTuH
vq+BAZCS9TCWL3HzJcOy167R1h2TgoF7jk+tiE4MriX61y/VhULyIeBIo+ardyfSRiRBDnr5ko/8hSov8aXEm4PRXTDBwukULs/saxUPkzgzLMvS4ZGvkLpI49lTy0co
SgWzhSZvGJq23u0R6u6usjodzowSrmQhYi8TNl1JGm2PYPSDNALM9UW68/gVW/Xa7D6/l0ZGcgLt8Qatm/FEp5hbVrH+V2oF7WHFE17fuhuX+khv539KcmFYzJWHNNEw
8Dl3HMwZlgrM4hI3O4YfxE9e52NpgC/BN3itSRgP6wu2SKsixHpwvQb5F5NtbCqIs3mtzaMtu4aLQ8f/1oRJKXNIMhe4jE6dqHWxuNeX0FoFcclBQNbwOAVPb8ceAA62
hSbtXc622LY9kVWkEF494v8pAfTysznqirhPmeJprAiUDy7QNGVafltaqfzU+pZHP9WvTm4+R45cIpKrytG2RrdtzBZi8JxjMX7VqVxbJAQgDJm6l4BqAK/xM2JkPqDe
hOWRn1PS8z0Risd4imNW8m1oPIfhkzUr+6aPgvA45sTxCSy9+re9JRIn1tL4klwpscR2i6MoAfJirngcv2uA8M6VkhinZbx5Gkh4PpY36fYYB20YsHqMyEGxhGkmNIB+
onAvA9XU0HvNctHWT1jTjD1e2dL6xwSp4S94oe3wjdmdePkspCNxaiO3WrEFTWaSEJqqreM7wqdWWQDIkmwydgyfwdTnWPzuRebhToI6/p2TSnfYHXapFgjiVPsSqo3k
99QwZ+OEl3kTN9/uqNuTwvS7DOIqzwVosIno/oaUAk6Rm6M4UzmlAFf/GJKI0OIChn0hQ5DmqhDbpSrIFdppTLhwgW3TSqjamCDFO9BcApQxDmohG/tN5LnEi2LgbaKO
V0TJGW0+AbxtVDOKx0x/Dkx6KHOu+NzrmHPBspJKUTUjnXtRAL8eyhPwCwXbT7GgCTGtPkyyEAK+0TVWOJ8cgmy7Hu5Q4opo+B5EnaAFckwuF6seec4Oa4ThyHsEOVgH
pcgwpt/uj6GxQ4DD2ggl15+VmpqvhDjrNFzd1mWAAao3/StRUebSMRB+WSMJ2c8ysNANfXb/4KrEFkNH7bCGq2vViQIYVLtfYe28BavFPgsEXYGKr2kISIkLhwG0AdIX
R9gsLNJ2LgHLKcm965fMHyBoKUBh1LL7X912c85lxLBdFe1XikHCr6s7ggOSzOEns3mtzaMtu4aLQ8f/1oRJKaKCEhMd/x0QGUZizYKSdeyP+X9db5+rNx3d37bkMBJP
/RpFar/ysBEUF7Lb8G0oN7SQv0SQoWczReWyZ4gLrI3EkgZCVMP/Ou3FjduJy8lMtywmT1B1y/NGXvimnjY8UNfBj3DAqMO6XlTTC3QGp9//zJTnD7bjYWJKg+cNlRWY
R7YPIkTDFORHH/8dCDFNP4Dk3ATCKDJPIMQueap+kW0hE+CygyVJJt1YXkFk1CfRJGf5KXWeFIQ8cr+yOX87Ecr3S6FArkCWpAfkrh7gEZyyOwrgujpWxbW182FS7q8r
Uj4XxNAFi6BWhfX7sya93RPlsc2gZKPvisIO5Op6qa3FuBJh+RnUAXkg8QhQn82Wbb+Ajiw5wuJiM+mZpxFOTl65QGkBwWhn4KtyYvhgz1nArLUwrqfEas8XSQErHwdN
RV6rvp7T4wuyhFZroaUNOQ2rHXV3UOYT7kOT2VsC/MGBTGiWFNLgTl8iI3EUdVJyiM/jcwI4JfoYMUG5x/DHVJKL5B45UEdKTX34WYxfaLGEe526nxRDSAfHYYqLhxUi
TP66v5r+UDepwND4viST3R9hVLCK2wWrYjeqM+SRAekkcQlw4GZAl8LS2XQAECXiqZfFmw7y+6a0YlNHDvos9UbyTC5qDzjt7LnvJnFS1jTKUVdF7EavIBNjKclR3rJH
tcSyyiRWwoFF6dhsUh/Fv7cmcMGKcq+VdFm1OmUmFbujaBxNGP7cZqgrLCpYrmbs0C5tEtdshh+RGTILSji78seBG0hUoHdmFHoYK/wG/wmulMOgAYhNhNo2IYVaoDYh
rEV4oWo7UtCrNgYwhhG/0+PHWesUHWa4V5nTXuI/a1TBbl/lgZZ5tuKoXbhcNCn7c+V2Po38AsxNzbtkYFHoUaDk8AxSh6ZbXgwmGnc02rJFkmngcOQM88TitHqJ6MIc
0UFzxwfhSMBrbayzDd6cEbnr31e6F2F4POCufUmy553Dl/mrY8wGbblcLDc4tPZJMOXpDePdNa+WHKQz5zPkL9vHVJRNsCWXujJg33zsiLoB7ReHiGSjMdwM3IO6IsNG
yjxPCVhqJH5J8bRBj09+roufKnMvD8FnjC07t0m/bsQL7asmsobBP+cm6jO2FXTSIhYKoLUeCEAvSvUQF94T3fxRlO7H1oNTJ/rMfB/Cdm7grVACrZkxJhEUmbMNTiwy
zgrlo6alXRZ50NpLVneIIPs0MwlpmNMGWiA5DHoh/iqiZPlI9otmoVBIWEO/XW2biYItyPi8AAfIlrTjzfDKWhLt9wCc7aCgEt+YsjENsPJ26uBeIXIL1nXIdouUR7LN
Abyvy37Cncd1TTSCKR6OiJPLRwTle9rD+7QJR9XHqLW0RtpnIB8AfcjVMIRqIBn3s5IOM9IyUozM4/OvDwkh6PCr4IGHEWnhxhKbnKDG9+OHdqefc6CBE87KOfRLZdB5
tSovNuaCoOL6OwVwaaZPo41dHMAo3ZUTV5//7vU18Eff+BP2d4FR1J65GmhZl1klxnwn7cU7ggg4H7z/Mz8Q1r07kl8FECSe3Zpw42+qK5YpqNDD0JL96pdZSMgidT1A
qxMMcwE2AI6Tt3zVJjLpXavGIDaBIrqYv4FTJbixRgSxNUlXLCaihkKawxMYEvX+Zau59l6VfBVUpYkGFzgJKB45YZOJ0taMCnyU0jaAWAFbOUNQ1uc05rrV1UKTi9eS
NV/NBs30LuKjkhgYE8eglu5BP2FyISaCXvQ57UCWzaO7Bo6AW6Ueq5u4rCrEWr0SLVBlMSvPUjbP++xP4ZyC/2wj1KCXAQAVX3KeMWaiRUEGhxXD8g0uWlUjS5jfc1XM
bHL/NQZOrSCAh/tGruDadbM4vyYkuX2cwxvOlojqvUNVTMBEKJDn4Txp7ySZwZAFuMHxQ1wU3aPN1L07ON3TuowAmuFCyLp5F5l+N60wFbIBX3TwfvAv7fbp5+nfgeSl
Yl1YuHh/zCmMB1AApL3L8bxrxCqzy+vpOJUfiVFpfvXWz7gquYoxKA3twe1o1NIhdQ0gDNFKi0rsOn9r1Uyk9FpCYidLQK/4EtODNrAx6dfCTnUPwgrsZUdVOMaxKGYJ
LA2nZGE8alIt7xqnC+3Fa6EwgckrMt5CIeWgQow7p2Df55M5sLATod0uhn5wcc6LXmOSgahwP7Ph0FxF9kffLbQa14Vr1s9zoN2b7DH6C545Mv6ZiHFvNv7U2AyOuH34
+UzMxb2tCZ7nVGRRVIVIYPh139E40hr37UY2yZSu2p3TFJnPv9o+UdwLAJ4Bqj+s8GpUAMiCGkIA2riPYON5VwpoS9JHdiqf1JXuzzvp+lu5CiaW4XZ4m023IUaPJfWo
EkLTmnFcN1lL4zAp5vxW/I/E4vhfWeTrdzF0HXiSc9PjnwxNnqqZ9VgUvh1/crtySNo2WuzA0AP8c4nBtjVyJZTZFqC/PXWOSP00sfWfso7KNItlp2J4io2prUsCONqf
keIAPSUcA8beaC0K+/o6Aea3XNUb+9ju/1iBr1YrQ9CNXRzAKN2VE1ef/+71NfBHm6Pq193l1gyYuD/nAU5NqiDKhbJbuqa2wCoFZoZERDN32vOjTHAZB+sZi5L2Lxiq
7Qc4L4ny3fQ/FtQ6XJKa0HWMgs1G8WRpcEj62NXyysuR2tEZQ7sAoJULif3TPGC5tVaB6bFqzPIlAHl+vWKLs0ad67fZQAdoIr/f6FvVALXZCSXuso0KtIKiAHmztXAI
2VBcSVC68+aY+qgCBLx5VBZjhOCZDPoCUaU+3B4+PcJFHsAHnOdPs5UxaiCYZKtWaVpEvbHUFJYt+f/T6cBXIPgLA3kUtMNZDXfjj2iilkABxXZvlpBuQIeFIXdfkRrR
amM4ojQZzbZPVPIS5R/tg4WT9BzeoZnXCWLzHho9ZuKoxlmZ+Q3eL08PkbDlYBjZvbKW4dhtD8SLpLB9bBzxikHW5lu2eFDDZJBIlidz+ZKPdcRpXG7iylw3JRevDFHC
r7pBFIqB+lfW564yIOFr/A==
`pragma protect end_protected
