//=======================================================================================================
// Copyright (c) 2012 Capital-micro, Inc.(Beijing)  All rights reserved.
//
// Capital-micro, Inc.(Beijing) Confidential.
//
// No part of this code may be reproduced, distributed, transmitted,
// transcribed, stored in a retrieval system, or translated into any
// human or computer language, in any form or by any means, electronic,
// mechanical, magnetic, manual, or otherwise, without the express
// written permission of Capital-micro, Inc.
//
//=======================================================================================================
// Module Description: 
//   The top module of I2C IP
//=======================================================================================================
// Revision History :
//     V1.0   2013-01-15  FPGA IP Grp, preliminary
//     V2.0   2014-04-30  FPGA IP Grp, support apb interface on M7
//                                     support emif interface on M5
//                                     support FPGA interface on HR3
//=======================================================================================================
module hme_apb_i2c_top
(
 clk,
 bclk, 
 rst_n,
 
//APB I/F
 penable,
 pwrite,
 pwdata,
 prdata,
 paddr,
 psel,

 irq,  

 scli,
 sdai,
 sclo,
 sdao 
);


 input   clk;
 input   bclk;
 input   rst_n;
 
//apb
input           penable;                // strobe signal
input           pwrite;                 // write enable
input   [31:0]  pwdata;                 // write data bus
output  [31:0]  prdata;                 // write data bus
//leda NTL_CON37 off
//LMD: Signal/Net must read from the input port in module
//LJ : paddr[1:0] is used to select byte enable signal.
//     IN APB_DATA_WIDTH=32 configuration, all four bytes of a 32 bit
//     register is enabled. Hence the LSB two bits are not used in this configuration.
input  [31:0]  paddr;                  // address bus
//leda NTL_CON37 on
input          psel;                   // APB peripheral
                                                              // select
 //Interface
 output       irq;  
 
 //IIC interface
 input        scli;
 input        sdai;
 output       sclo;
 output       sdao;

//protect_encode_begin
`pragma protect begin_protected
`pragma protect version=4
`pragma protect vendor="Hercules Microelectronics"
`pragma protect email="supports@hercules-micro.com"
`pragma protect data_method="AES128-CBC"
`pragma protect data_encode="Base64"
`pragma protect key_method="RSA"
`pragma protect key_encode="Base64"
`pragma protect data_line_size=96
`pragma protect key_block
oSWVujNS9cA3DdfENxE05T5gcLdoAZK1ZM/dq4NBqboq2J6r7Xz4UA7p6IeIGt9LKnXtgwvfhK6hi+sVIWNihGbEAzFSDPxsM++Dr0gN+kp7ZSe1ly1lBKK7w8cYxKQGiFAVX5QIZUmaCrCV8eaEw3MqdFahr6byi8gZQhC19bM=
`pragma protect data_block
KODZW0d0VCrsXIgzugfefU46f83jLeI09zQQUoU0HWoNVtSGIkR1ocTjF7FQYAr0KODZW0d0VCrsXIgzugfefYwV5k6jmOXCIJBiY1J0LDFPcyYJ0YCMdPROL7ELY0l0
RwZkiJbDjpThiSH/zh/aY0AdxBhcusVJxCkdNDOZa21OYjFaKLSTBRuSSsLzKTcWEgbzBECOcmhvfgnS6t/dViCER0zi+Z5upVUczL17O6DQUz6QylzqSnEwKKlcOM41
FCNIRr/QD1L1KmNeAFWvvnXn/+i4p/w7TJ6FuREXhPC/ytGWxwLzJT8+TaKV+9KEReTxmicb/N+ZjruRgeG2nZA905hqrbnYAj+psBmRvnDGvQP7wwakNGdEww8jOqHY
OFp8l7u3iKvscA8Gvbz4VBdNP3z4ek4j9EQkwUCNeKa44wubkUwpV2RoWV+OHQOI4RWpdQKCyIpcz7xSkZyaxS0ibcK1p25nU3tK7IJcQ2hj0a1RjWdDX3y0BbGTHFee
32bl6et84LWBI/q/izTrV/9eb7hwREf0apFpzw/fz/n+nx+k+Okp3LJNc8NQ6lLVSKUEw9rYgLkrI603kr2SW1fI8gacvnR73sYOXlDtRq77NqMyK8J5AZ3SEPvI5FXo
X6PbdUe82yDOVQNykZaClqwpqix7Kkkxx7bjm3ZPhqFuXnURjpNE7APb0gnrr7CuCIN6y3zWnI5JBDSngbmVaduOcGvKXlB6e7KoBzITauHthuLRWKfFjlYRv3hZwm8W
LXQo8l5EINm15enrlbl6pLqI3aXm3tvPX79Qymj+MtA6t7mZmRFDGMX7gmjyKSGSYQBU1V9osGkgNoC1orE/cdrNZ/7p6tyDiFT5r2vj/LnczUDP+Kt0Jeai/UKYrmdp
fsFqqG8FfCX43hHlc3OzmYmLk1YI7S+PfY0hmlU+XAkenFYnGxRJslyHAupLZJlwdKX/waO4RciZoDcbE9kr8xZPO8quUs5ldIVezxYfSG1iqwMB20mNOXjevaQqcLp1
Ix832tQDGXmqaUoaNXw36Dr1QIr2PPRSci+HeZKhuXh3BTR6N7JI7puAxpwbNV1U05UyiORajOs3oA514lgMhTaNILbABmaIb3TXxpbKGMdRvuh/VsyIza8KuFgtG/hM
jvLd0krzXUFhJ8D+B6Qpxk2pza6LznLV4lmOR9uj3NmQhSJpLKzQOb6FFgNFnm9v/JivR7EGOz0gKpI8Qu5n1+gZvktOw+IkNFoASgjXft5qk0Q9JyUg0FXZW0UZa1KQ
LArrBQixhhHlRcqs1DmAz0/Z9t72lskFGChcQE926On1lE9yM0xzsRG6rhMZkf6x5MmA6ZhhDewJwOdxMzS8i/Rl7Y+Yi5vRVucvKaHSSqvvTo/6StLdKOUYW4NQzKX+
xhGzFJkzrvU1WAhoD1DxqsPB645Dgs+5tlCQ5oqBwhZYy6++dKvtVmKmJwdpfqtUeYv17/zRSwLBQ41xNIvvr4e15hBlIKgb5FWRLXOVEtrHG/978tWoh7hrrorcF17X
GmTaRqCVpL8F16zRYWNt4gDcGSN2kJcy9GR2dB5JwXbJtk0GNO9Xy+PVs4pklwnB7E+pkKUvYwu0OCbJ7XPitC6PIGWv6V0JHbGynOkaY44GL7LiajoOoZL16Q0Ugyjb
n7/F3UjmUaBfzS6olxz1SmjjP/lcqLRAZh5LU1Az6Oz8DdKmexq7ibeVTcGO30GIHwNs1gLUQdvgKxrQJVQ4Mo0YU6XH6eg0DamL6nKG5Dtb1KxvCt0QISdYVUpPJ5M0
j+ojbfO6cE8QS/LC4VG6mu5gZagCjtZt9U+MWb3LmZGc6OVYcuV310e7xKzgC7Wujiqr6lA/DsGWZzwk6HmxeXgFdxfPpgvvLoQhhIPfG90PWLpWCdd5iS+QdrErg0/A
MYvPleF2LdhiTRfmERHQLrk8Mi+1DfiOwSiZlq6w2FQXB8Jjf+R7HZ0yTaw28wahDW7JP/ZKIxo3/U4gO9jEpbi+DypZo+tXW7j81VA5c3qOF1/mbFKMM14xgankbVua
DMnUYlMasa56P5t+fF6Jv6CXwCdXq9KAGY7dRhbUO7VHhbVxwjCzeE0xyeQabm2Sa2hexPqEwYQvj4c3WXYMHESRuGKazajzbz/HwuEvZJYy8j7a/tv4MBmK3xl8iXHy
38uRnMHXLTcv4oX+dq836kSRuGKazajzbz/HwuEvZJZFb/gJKIfewfkei33CnV37Yrw9W2tPjlYq6gUbiOSo5uleqEZLOULWBe4SA+YYMg3n1vd/B2IpzJ18WWHfYVPk
XjQMDvRf4gq6R+xGpvQAtgSzl/1blegetfy3YxjLaKvKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiDQGoUt5IkEL3EcbX8f6F9we1jbRGIQxTEJ0UgDyNPze
EIeEoiiPyDbp9VsllxPcwPYYeFmtkTRZw6dKCM3xZmMBUzkwLed94E8POOLbNMuRyOYZW4EQw81bbip6Oe86rYS4Lny8fI9hR4rSg/No2ylCYlKysnbNRQ8XUgCQ2fGp
qq265vHHvzKN20/qLENWMECLn2ltOBZtdbGH3XxaDXk+ghC8TVfn0VthFTs8oRPEF0sJLL9wITp+Pq7qFXGg+hXtu9m3oWciJyKo4voCFzLeN2bVShNGnDxzzPpyPSNL
94eehzzFicHAzK6t7v6avFjXacrnaLT4HNdKY3fBjJuO6PqvLeQAeYfzRAhB91eOCdICQsL9O83+gqkwE48pTjGx55BJjqPPoW35H6rbqZdBxvd0G4+6Bi4Frp45unj9
YrM2YFVH9gjHw8myfpxGzO1QGjM6jBNEff8VV6kZiPRikGXjJ85H+jfgW1BAVPlEFGzof0K3QeAIR0sNbHA5yoPSeLNp3Ocg1SUCGsTJw+Pqr3yll7MRZNsPilhnooPk
KkHTYLZ3eFVgR6Fcq8b8rAwtyVxHvTfG50Z+/45gntKxWtCTf8kXJMH6bi2jMKq4dpK2/r7L98nr0zVqnySGXv0INw8zixlGlPCLQhKEWgWEbAoaFs1UV4GQftX4cbz0
v5j8FBlPnD8OE2eg3D7Vs1GVS9CEwTUzmiYZ9DQH01aWOHu629k1WbHklxB+O8zGuGj6T8qUN8E7mjca5YpwTx48QI/uwly2PdbX3DwYkExP4AeQV2BWrBSPnOneOgWS
Xqm7GfrJXerdSkAPbkTOlKaRAr8n1d+O3gAWzvaxAduvKsrrDpfFP/PATWZG1z3nnpOc+s4kL00I0R82wyjU3aO0nABY4/zJvPRkzSNyXeRaP0fk7dYS+QUJ6cCV7r0/
YfQyDv1alSmnKb+vjhcIf+ixhNiWrwV34SDQ4OGHvPxdINdIxFXF9d7W/H5Y5lDRLiOSRUkO1aY58iWlqqgb6mmGtSeUZyrV74q7vgO++NdMOl7uDZYRzqMaCgSHPArh
Oht4CgrLpEzJXBDNTAXmrDrJNKdL6pAN0UCSNjWEqTv9IrzpecxdvCjL+2KnDjbKJwTfuLMLvu2KRs7g/uA2nZ1eYTlH4d/Te6B0W0VG4Un9tUkcx6PpopyOa+s2y0D7
CGAg46kJPC/lcVaH2BKcsJ7dTBo8kQ/mST5EWKzz51Xqr3yll7MRZNsPilhnooPkBKCAcS++dZLh4zqsjRWFHPsl6cRPkAtL0dZ5iM2lMS9huNDXxhAaWeQpPNzsxeDy
BHxMh80eI8BQwG9kFfubDqrl0g9dOXX/PnTOokh+fSk9P8ryCL75Tdh5jkhK4VgF6c/0RnpfYO1QyLLFkpFDOJElgCOEajZsMeYkxm09VriJ4v7JgFDEkD7UfPEeoI37
leTWQ0aJpgJdPtfzDRnV4ugqFhRnm86JpC7iFvyE85+gJ4aznELqy0vexHQVv4vbpjrCG0PioY/uB1VaMVovEwBTn/7usSKbhfxdKPXYvfgA68/4j+FZgx89R8t7L9rg
hJGEQz+T0K9AniccVVWKohPqyef+8Gr66vZBPV7HoXyuyuX/qkuCCem6QzkY/bfdYxqJChXzPl4I+xr3YMbQNqE+iMpSeJICAObaHfFHk+87ZsoV2xZ8xc/zDoi/zlfT
sXgKqVeNpWeaq7e2diBfVN4B2DQMDQBXDblvIrWw+tOJ/1h9eWlqAYPZzhlOryV2uar/LV1fKDVti+hfP2A/sIT2Lq5Aj4lB4KoP5rqt5SSMEGEzZv/yPIl68fUVev2I
+rBHuSdI7TqHV8vyT63ekjatJNv6hY2DIrY6C6mqRlu3yevFtwMmz4UI+MxG2iMhcCAGfLmPa1thOWVv5dmgC3B9mFxW4pfFwLU9230hwiGmuCAd6+LmrlBmiFI0EqLS
XDH7a/1SMrnJL+kjz+BbP8McxJmPbGcQ/tItpv8/SEO/JYhkIYI/75ziBhpjNqsP3PSu1P4d9zAvdOSn4rixYQg1ZP3m55izMqkb8wL1JBmMII9w8F7ZFsHj5mb7t/45
SeqW56pYxoF6V+zDjROISfJjjMNgB5Qf1gQYs3lsKwr3JUKkOLbKqpBTI41AKYy2iIVBKUPDdD4AEK6Wm2dulXHVCCLo4At4VYXrVginlYqtR9B12hCsTW1EF414zMNJ
cQHDxseuKJ+0UleyyUgfcoo84auBDcfoWrtY4tJxfc2OqDZtzaWdHunrlHrgMqhRcowo68W3qd0LQmfvN9x/Rvaj/Fo4iC+jMJGNuv2rXPbebF6p7DERHHo3ck6PIBY1
sRXHdKkLkLePBUNO5mi3hwR/PB3Nx50H0Y7FsAn2hN2zGB5eeGimCFIF8CikZyaMiw2uA+w+r8g/TCK0NXen2LJ4PLaGLeNrP64Y9colr2MTqY56x+1gW9/syfrXmObI
xzSlbFOi9w/E1h7Au+9bSY+3RhmvPCQuKgGDdBjK7UY3RAvt6Z+wCEyr+D4+kGJ1Qie0kEADKEjbBDqqEIPIKqe31plynCcLewsWAtQamisJZz0BFgmEV0FbWi/MQ69H
auMY6VccqCsoV5vuq1Sf4EoJ2HD3iDqd/nXyMTM1tNP7709rDAPRbtLwxtypOIEh5UrM5hS4t+HmOFE4S0+OBpINimGbR0GmM16OKRuoJjev7slPmTofue0D6MaKf+FL
1HfLdIkL6vXvk1Iu0vjcW7WOEKGOiVimziY6gty9oeRsHw+ZHvd50D7t32cSCp92c4w0317lFOL/eqDO2AOA21Y1JHGSbF7kWSH9SRHDKrePpLmVtm/GdRrHLCJhZOYz
FjffB7yJ4mYQXq4h1JaafqK5ZhrnHaTAAtW/UyBlwDbSb6AVacAWRSfxvBpmwtT7d/+LY08PwWSKk2o1ei+clbv5x21lY21uy56amT/zNmKJSBkWTJKHfymhSTRYY1Mg
fDFxASvq3vf6UKvB5iIGrNt5dSkH6OPs+xOe6REAqmc5uqYgKbZf9do+njnZ7vscJbRIW5EucNAMJ4woaQ6sYS2jT+AX0hpgUD21VNZL8EoW880cZUmuWJLKby5GFAPY
TpD3OEeoEahHyKQbJjr5ubgYyBMxpGZK+z3s5U9rxqKCqS+PB3RN3j1wfzXIVQPinQx/rGeNdUH5bzNTgazu/nwxcQEr6t73+lCrweYiBqzz6cwZMLwdBR5NkgL98UUT
JW5joSGxJJPQu06gQnImcE1/dFQI+bNoTdA3CtXKYvSWxQEh+Y3lrUeC+eO1rkewjsKFsMl7zqdXfiJdl+Yk4cipD3lQR67zGm2eipIkgs6Flc9nLF4seoy1yxz+IXZo
Tza+RTbxNGt1YpkqS40/sObv645Uy/3s9tCcy3EIJrTq4ktinIoa+M+J2a3lovWd0Ubrcd/0EcDFltMQOcI6Rd3DpWLNFn+3Sc3/6aMZWff8i+1QHHSsGmcNeMRj+/VZ
wBz6WHX12bg7k53XCn5NJWKuwKyC+up4w7io4a4w2rIgZxuHLatd5jh9KKUnwrnIaTRL6lXawyRT0aEAvMw/Ntn1PuUcm0rXOYcl8TbCC56W/J5hfsfyTjI86qf9MUMW
7saci1Od++5P3zCbRJvOVgheOvlkPgMsprU7NosMddVw9R6MGklTukDaxHCcA2ixKT/KcCXBslhXRHzff5qHgmfk5ome6R47hK9LhKvhEuZEqg93J4kyHg5mskW7Y0Nu
WrYrl/YOeyxp2pOkvd38DQfqd0vs8XOuoW3mjhdBdqb7YQhaSII79JJHSi9cad/f9b5vr+IUeSSvtMPS2VFgpp0J3152GW76rZoD7OWowcskL2KcY/D+bfeNCSlB5UuL
enqKBMHiNz3dmpMx655B9mbd1vCUTy/whIMpqNvMRyhEqg93J4kyHg5mskW7Y0NugAr+6Ec9OMcexeBSLziZvAfqd0vs8XOuoW3mjhdBdqar5GJQDMcQ1Hdk/Pv1RT2N
9b5vr+IUeSSvtMPS2VFgpr3JM1ueS0sH06oSz4q2upVxqNEnFjddp6ted3on2r44l4SCKQTtyM5fvMdpfMXafZyxjjWJrrwoUpl9kiixdcoH6ndL7PFzrqFt5o4XQXam
gK8SdZ92OLTn7q/uYnlDwWm7Jh3pJloKjIC9SX1CyBXnyXgG2x/LzKVTdjAf6b/xlNShphgC6XUTMr7lHfaCakSCsjM4HIUACpK8332BxrbdodQpY7n812nCFLm1Chkx
iMHEdFrFm/RgLlomDSGAdFtQJQEcn35Z2eoM9km95+oTMXFvhI9Pd4eoGMgxAkolt/dzoCtrVmggBnqr0F2+gWbd1vCUTy/whIMpqNvMRyhEqg93J4kyHg5mskW7Y0Nu
+HLnVf/6ErXR2ZIv8cEVGQl5/QP+s9Cq3KlPIhnCwUWz3OWQ0GTAYMg1AHtcqNJeWiCGe3S1IOEJZOeu8QdokBxytOStrpE4rbUHhzHC2M7tHwY2Iq4wImAH6ysG4Lov
yZ+Y4Y4VCU9MjUz2JpyVsWtR9o+9s5qiOZdgnKwR/5KqX3uZ4XktStFi3wMP7A/UTsz4FJDg3zeTyjjDpItGs8Cbx5gluwBfEcx9qhrqwDqyx8naRtqjUJzMx7bUEvSr
Yo3mDtr5CzDiRcVSXnPMngl5/QP+s9Cq3KlPIhnCwUUKndUpz0Cuol5T9zm73Vf3ARWsnlXZNniN7qDztfQerKLJ1+gWa0rDo29O2hmbM3jvcL4DuBxBOoQS/aqixbTW
24wdCMnQWMwuGGezr0atBUz6Yn5oVSNIWg+6Q8t/iIyMi6Z/hJ3GYRXCg1a4qKXMjYAlZzlkf33rPKg8Tkrowbcy1QANw7ARqkMJIFWZNs9EgrIzOByFAAqSvN99gca2
jnTO9unOCxENmmOJ4rHh+p6TdIE6jmtXMwRCIXb/o4MGriqQLNxzyD4BPm+R8/BuEidoIy6ESkmbMhzrQS3YlMmfmOGOFQlPTI1M9iaclbEGNwJQOjgZmVcLYm1kTxbA
iMHEdFrFm/RgLlomDSGAdPwm/ovIDIFOtNfK/qSTAC6AruACVlPi9PmdQSdj+VIJSpc3oi2kxe+/S/nIJ8U8HsyQvkXOIUNoEwTJb/5fYq4H6ndL7PFzrqFt5o4XQXam
gCUuJa/q0fz3xs3jSQG841larjylGu4mU1M3VvukWPSXQUXPz1YXzyjuBDed0rkQrfk3cLFnFwFVMcmPYg6xEksKeL7VG5fQIog5f3/dyyLuDPO7THdjQsVGxfy43K97
49ga31UzPDP1vJXCsS+b60hAxIHZgz4q5UstnmgH3ERuwUh60vuN8MrO1E/q4xbKRKoPdyeJMh4OZrJFu2NDbhppQ4OWX4ErcBLBLiaeiKk4elEQVklekLGdvDlUlSec
Bg3rfD5NiPlNDlkU5zw+WR4e6h4RsfeyZg6Kyv7HKC6yx8naRtqjUJzMx7bUEvSrZH3umjAEY+ukaUA1opdb1wl5/QP+s9Cq3KlPIhnCwUXrDG962B7GbxBinDFQ6VG9
6S+ESfHLPaTgED1VyZBwtaLJ1+gWa0rDo29O2hmbM3iWgFIYPgOt7JlkQ/9lgBVP24wdCMnQWMwuGGezr0atBSEjz2i7Q/aPwquKH++cqzSMi6Z/hJ3GYRXCg1a4qKXM
xfDGVlv7KRqTE2ZWzLxs7xS4RLhpKMhmo+y03QLxen5EgrIzOByFAAqSvN99gca2WIhJoZYNnHSmHDMzKoL5tZ6TdIE6jmtXMwRCIXb/o4Pci4Lesk8qPywwen2qWCKc
el/wEef10zVJyEWaHDUDUsmfmOGOFQlPTI1M9iaclbFuR1my8+SD6SnUNSHHa9YKiMHEdFrFm/RgLlomDSGAdEmEu3qOdKaOog9p2NE0HyRm66QiIXoHREdBC8jeZ1ue
Spc3oi2kxe+/S/nIJ8U8Hjo95CzW3TIDNM3//hexehoHAvVgLUaBv210sKAgE5Vvnga6yN0MhWGcaY7ZAdmNPSlbZfB6QuW4pw+S1Df6i0NMFOF8SKSOteePaYXk/Xwf
vFfomDbVGSsZ8Wa+5LEwvswVVUGroHjEUcyeGwbcYC4h0e7ABCOYB7Kv5LE5np/iRzdW2YzfuDPPjzHDWonaY17Fb0KkwhsjI3J8/W2SyvKIsp576oEfaCNzHf7r9fNW
tpIb95n66Dvfkv7NfZk934jc/jnHlUc9XDOxnYpdRAKyNjVPlh/bVTymXlqZB5jXxWg3+pa8PuIql8ufWqFkod/pELnWpnW7vT7c9fZFXfK4KQg1MNXhgoY5gDJSMwfD
6CSxxUr5ZNWhvrdqDZEe1TDaPqZxQTawy20CnmJQJaoAj8VCvFVgCOp5ooL9X1YWfrutkO4SlAoLSN1na8GxrMeKEF+N+XNLsS1vjaLb8SDnZC65SgfPC03+Ay8C0u3x
RE7SMNPd5kOSVN24V78w3mm3Z2oUvmE4RTEA8aYXGrW7wkmNQWVTPPat9VEFfs8oM170bNA0XqWJz7vh75yc1YQ/1OAC30fR4BYEs6QNbAQYhtU/I0trNrMXj8xfpRo2
1jfAhDMKHw9Jgn2I4LRCmphOd+ONVnpcCiWWADL0ueM659+6UQC1ELygMo/fvvJVwo96gJZOQ7NVCCLRFGkq1hAMd06eXej5BDq5xe2yWS8oMOVGIx/yuEvjhk6Lxd0P
SsZBcA5410QXPq56k1VH6O1g7vtTs8Cg2oab+6sDSEKioQTzgTnxugTo0vQidW5NxPswrV6BccawJ39O27hFU999HRH5M8Tie+phAG5Ke8Aej1ra6XGW9ZTa+psNqtLa
XEhDJ0jyC0dAlvPPClfWxDSkdVvlpHa9FSYGbjQNzxZE+AfC+3fWukAM93VtAOCvb15j1/luuMqBjuQKwleNDNieue1NPu65srFFQRqf/e7oU3BlSdanfmgyyJI6o+eh
sSlOJB6y+fj3WyNmn4AWeP41gUxjMjoAAfHSQHv4qJJBq6qYb9n9nnSYEuqXjC7WZGObHKQJlMjUR0g92KIDUyAC6VsdF33tBM5+pRwspwPZlwzwiaaN9Epq1IbiZ2Jo
yUE9BOzsozBCfJ3ES6tuPXrHPwn5R5rZcsuPytKmlpHe5uuOb/1sDSqO3vwOJ6pB55O6wy5qDOTrBFG8sP+MkCKUpqi1YJkblF6FazCDI9n33Je4du6muBaHjJBDjmnp
XoiybE/Pp8AZvtpgqpemBSgw5UYjH/K4S+OGTovF3Q8sXn1vGjW0LYpF1cCGgansrA8yEGhAsF91n/FxwjSS/Ej/bkR6fQ5fJ53gan3klO4AhlWy5VZfCHp0zPp7qKYu
u8JJjUFlUzz2rfVRBX7PKBlFa45v4SpccO6oE2lXH2jl34ImbPhGopyfip8j0E5o4Z8/JybzRV5JC9+6ZHbwcOSDnV/Eurhd3+Ffz7abLWViS6q7WTZXpais7UPvr4Lq
L0aOYQis/1aok+iwV1ks+CLnIg3NwJHb9+iFtkHm4YhrRg/9e61/0SRxnalOTaZh3ubrjm/9bA0qjt78DieqQeeTusMuagzk6wRRvLD/jJBaaqFxrpFG2EkRnIeaGoS1
HpQEcrYdBPxCeU3OLilvBTxdBXsN8fLfnBmNzs3bF+dJ9hSISZnKY3jOT2GuAuNedbbZbbkfv3wJPwDJnjGhvClH0RdQ7ykZukL8EjBeubrKLPEn2LavSmEZGN3m1uy9
WECAHJjRlNHceYLPqb8iFg+WZvM+9kkEj7t1R5OSO7Oe6yYmDJRO1thYxYUMC2gsp/oumF0n8r6mi9SgqNT4Nc8XAIE5ryhNoe/y4TXAMvseH2m84IJ5cy9yjYS1isyB
89tT+ydKbspcIJ7OYqfVa6Nl5PynHMBUXvB9RyzQg1DlzERm1//Ist/QfVNeWL3S85i+HZePdWA3Ocd/yEghV2HR6lDFUepi3X5UcXYvLCjz21P7J0puylwgns5ip9Vr
08yxBI6gvBZJNJU+WD/2HURGOTvbzzaiVf06jH1S+h6/iJ0UeCja265qSCW3a6AM/MUnb4dzyavfn1vUMJvRScWWYQ/NrqIgxduaC8QgwF7n9ZpieTmxJPcFtmS89EcX
hpc4iarZzgui2KCbMZhWETfFCelgph8cbixoTNXer358b0mvU65b0poMAYPskB2QRKoPdyeJMh4OZrJFu2NDbrfJplR70QgA52FS8KM6a1UH6ndL7PFzrqFt5o4XQXam
BEgNNOGjJmJPrbeAQbShVkgeUD7BfjMhVrei6dcKyUqH5UQ8BENSOrWSsM+qq5BVxZoT6QIwcTqFwnIcxPPEITfFCelgph8cbixoTNXer36Ry7V0bLdTjN42F7vH16+I
RKoPdyeJMh4OZrJFu2NDbsk2BtzUdMMX8/bsFiEbBaRr3kIIOTYM+9EzeNvF2Jai+tF0lBh1DARhC+9GK9A42rntEzUSMHFxH3NFQTFuj1XKiCbRJr2HgYyrX3ljAm2I
YHqOYjXlZ0YdCQQaTApyQOMR/5/rORpcAptc0trQxl3hiPbVKLKPr/E6p7VmCPRKyogm0Sa9h4GMq195YwJtiBWjkJBTCWJ3vXqnLrw4/SML7iIfq/BDoBiYqO57Fbp6
KubFwyDhLTK9NoGgxbq2HTwxCgWD1KOcIJXP3V8ErtOSV5RtLiiRKDaP380zyYneOEGmQDr7FVvpJP3TmFP5XyMpnacqJ90pLICD7f2zhDNNsP0Y/DIZx1NvHguRotk4
EH/aqWNSV/HGCd2MVNI/IzhBpkA6+xVb6ST905hT+V8BMn+9xF+QJn6B6uhwcy2Fm7mMdGaqT1tKEbGimMxlglvXxWiZuZFWJ/U9eN5jMmK2BUqHViil/f2QrDLCbFX9
UoP7+BLCznWUvknd5/N6hCuyXBsTzbYUddvxo3NHHDAlV+rBKcgXYO85M6yWNcywA0igMilXfyLzexvvHpIeD9zUOFWVbXPitQ12zBukYhlmfZDuytXCrQ8Geix8wiQB
4gGa+0feTza3DJ4DeXP0MsE3Z6KlVFhO0Nd0orPiYYH1rtc63sBvoIV0s7plEYfekXJ8vXvxTjhIT9K0dySLY77u+U2ZGOjLnBLBi7U9GsdUHVIQFaNu7TzPHmDAi4OR
7W3DY7V3XRpbiUSqMlXZxWUClah+NvLXyvhm82zoY99XjJnCM7g6MnqLEn7UUGi0wz9zogC4MSo3wD0OAEWjkKR52Hq5ObmSizNRkp71KlcMXNHYuZ2ym2MpuCAXvAvY
8ChwZ1oXqe47MYQzxujXraGO0Feb31LJ5hjl+vLv8JdmfZDuytXCrQ8Geix8wiQBoZbbzCtjMvHElwgZdXOWVhEG72KXvbTgA/xBi3HXFInbdnvPGjbam8qeNQxS+sI0
CeZh1Y6YTTN/auYFU7RRzbF+34AFwHDkujI1VrAmXpq2BUqHViil/f2QrDLCbFX9ESyRWgJYqXnh3mJKs8/HRfaInDlfs7L29133xI5onuUtf03UMUBGsWVDuhJiVRAC
BEO/ApSdhbAXS/glpeguPcyJ4H5w/xR7gQSLW+CjWKwOJJkNWr73ntwNP6MSL00nm0OcHdvyivtXTN/BROoxWkjMXxySylHB3cTbVsSU1q13u+u5DqgEaIgCJBNXfPCc
h+j+ui2k6hJZYH+U33tUJu7uz58dnxj/krxY0GM3BMk5dRXVlTyGtrNJI8eqJ9fuGruyWOyQpwyBuGIDsC9X0XR79AJS+mZ8X9vx3Hj1bQXHdlAsquXrFq1+39rLQfR2
oKwGFpH1g0DPuD91EaIovY+2N7ie+bMMiz/sUyE2LYfVpeVaWkNsGnk8F3EUiR9yWigVkQwbuDVrNSow35+PrbCwbxT1vDGtGs/cDVqT2bPGJxoySZrVU3COvUtQ5NxO
IzYGf0Dxi0cN9ZPNzDOwgyG6o/6bBfIgFkTyF4BCiZDokZG6pc5LidvG4Z8ur87ObSz/gqzYuwQTg19u3bFqYLWo8hhS0kHalaH45UBHnkBbd0KjXanPUh3M9WWITvl5
mgTr8Ro+hVQE3tIi0x072GtpXKwRsIbbx8D+w3ZRSfNJ1TxxfUyE8Qk/YxW/TtTKNvWZm1PgYwi7+iNkp78PTcv1nwI0v6Bsuysp22iMQJQWyEteLRfYWiVYimWmFDjG
SdU8cX1MhPEJP2MVv07UyrfMGyYmun+KhMHBGIfsheG9M8wYf9XeWe63KLNmVKGTP7iqqLM8ATBugydRwnrly76gU5AAGNUVtuJb/Q9h7X+PnOlQljoeWH3LNtrB6Tzt
4vRm+lNb+STFHtMmwEoUpjQyNY/aIm3uomZOh3/oxw8420YUgf1HXSMYBIS4uURQLozQKOX9I3MU+LFzELDQiKB4MVJg4V5PZ6/dM2XlTygUtpO6s92oad26MkdPQykN
DXBLxmpCzNNLAuPJnyEE1Xb2ziIMgphXqT8NBCh55+xVlsSsjJp/7SMG0oLZXbMygGhiGZXl/ol3n8GZ8FSUQnFVv5P7G2BmIVd9lIjKmJUZaNzziMgTDMa3NhSMC1Ez
LFB4rOMCadMe71ZHnsZxjVEkJHUm6YXswprr6RPl+kt29m78ySKH8kIYFG1RWXvBImAKptWll9modLw6o2KJkFaVplYUWkmSNImHaGbawySBBLoM28tBIML1E+WMBNj5
jvVfSXRhBkefeAtuQ7vUL/NolPFAlZb52uHZZBduWY25ZaUyZjr47W5/JKSR4X+IQT5t61O5TSvSmHHIz4cALeBOaXvFOFsRSFlHWbHPqvlQ8Bu1jDc6KaQw9rXETfaw
iu183B8wHl1B23b9GNS1E/1p9v5Lr1up3XJtOvhLvmSzLipTB+x22Q2UTMU1fM0qWSdswL+IDxzNN9yOUOp6ob9uuWpaE6z55l9715FDCnS8drBE8mBDcUV9u4IV8fu9
kK7yOfIZbszQ/MRoM7d+syjB45bpHUM4lW9Yc29yYoGPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCeMbBkGgok4bcDk6sa0jqR
edjS76GUDXn8KEgAuQSz2srY7eX/yT/l/TPWlRqLqeePtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMBaT7mYDgfA0Dh55AzCXVvh
39Oq4Zak3kpdnMLViqLh60hSSX0+mRrRufToY1RLKR+8IMhcdY7zSlNIE1GC0oFeGU5kNrxkQY+V1wbc4hY+C1OJ/dUptxVudqN+HWiU1qk3kI7LDgQh3dKUDmiPp4us
+HfzSpJl+TLcNaEat1EO8UzHHFT14SNQEpahaa7/6kMM074XjlcvrQC26AEzobe4wx2+4ykhujdgPokg48mf7cr8svTPkd+QkYRalr5BAnh/1DbHFDie9EU7tq1lTUAQ
t+PjlmS5WbWBQQVyKijWt0Y8iNVFULFqWD4dr7/IkTR51Kvf38Vue4RSOlykDuaiRBsz8ox8Wm4SOR9dKUd5aJO2ErpsektwcDH9X6uAarCTYOSOhhzyNmNfgun/pFti
fzo/FMSMJ87BtwCrut4MuI3KeP8MCzGR1kL9Mnb+rN+Bv36j09YaR6BI5RRvLEz6AFqWZm57RBjNodSGevKFKa4a5fuUby+OBD5jzFhTX9QAK9zMebT/6qilVMgoDBbh
u6o0MbqXqRanQNLFBxgavp5/7ni2mlDf2EV2/HSSSeT1RB+c7dBcFJZBqmDKuWpZxDAKKRYHmIow7A7dBD7lGZfXgsqwhQnu+bUNU+yaSaPN2kPwRKc6+krPRxQsYiCh
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAiRO0Pj4lAAl0iKwnTZNbjH/rqCdAn0+f2OHXDQiIMbQHiVcIde/tlZ/mOe31QrbS
Q7W6nagqCbeGw9KFVzU9556/WDE1EE0mlyyrDqcqzt2PtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMC3BLgSIr22jbN4gHBOjIjf
4IqZCQexYSwgs7oM2Tnck2F7t/KiCN1TldijC49MgEspQMzFdJs6rRieGTCECDa2W0by2ocnKsCI62hritvfFwnIkYJbTh73maaW/O2DTVwBnziDHcuPldEe8MD/0Zqz
9OsUJlK+kP7GJzlzXSSsfZS2P9UMv3bxS2Qu4eIcm0TFfM3LN1jvYOdorUc3wUfn5bEdHbg8Blpy6ozzmIGxD9ssE4/0/N3UAbqpQSPKqXdzjRHT2ymkRWLP5qVF94dZ
14EQ5oupQz2jeAkAkM/5tjfyLS9n07L+b1tPsQVH7ND6my7PnGd+eYlL5r32VDSGUFxgcq0FroYPPabyBClmIY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwJ6xVsOuQdDZDY7xXgoKe8ApSQnpnKNnk+6G1jL/7ZXGCknO6q/DAdTNWXPUCEuRwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwAiArwcu/dwGmi2K1BBfK9TOTqEPsPlp3yQff16Fkjv7ZoPfhm4vCGwjwjZLGzdOEhoj9nrN1IesbxEv6gfvhdwNdGqU5Ku/Yaup/lrd+rUG
FCKR0+Si9xTOPymoX9vfYFFkMWwQEPPaZFttJqTxAUel5f0ZE7yChSHxO6VHQ2QZyWcu3jRCr3DxKxISz3TtctaFVmoxJwCiqA+ZSm0sBGRPnVVeGeJ3FiRo07oc027o
JRX2AtiLz/RltWV42DrCditjPSp9hVhc0stSVS9fOy4WZiaB17hXKjIGSm8N82rOBbfGM75BnpXg/2N0xrSWiY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI8qeMp9yQj4gifY2gYG3nKqxWPk3thSygfdHnD7FmogVe9zBil0sEScg8BAcyQE/Y+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwG94KBrzB/EXi9Cz6+ft+hPGwdslUgrhNzLcYIiW+s5pa8D8IyfRtINP52vh+Gt+HCqefoJsgoXbO9JpOiiwS8uCZZ9rYIo2l+f4yKxvZ3R2
a8D8IyfRtINP52vh+Gt+HC04Ww5lj3QaOzwAKpWnGt7QvbQsnoYSX1ZjJHdECnswj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
kQDLA5KzPLMzcD+yhVPo2KK06lIZVSTdJbv1jTF5xosKSc7qr8MB1M1Zc9QIS5HAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
kaYu2JxZla0kY6a7DT9LoQawkAc73niSD35L4F94BcaRvE2KSnZln68RbcAXKm4Eb6t73Vb8nJVnn4yHCVfP/6qUcUoLIwlSZORabqPKJaRWls8DeiLVfZMeSFSktGr0
5I/bO6eWuV3jgnoHW1Msf4+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwBQoKfb+pJ1HSUdJo5KAsuWlUc8F/i8J5iH+urGO9/Vo
5RHAtCeQxS+x9mFcJ5/kzo+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwG94KBrzB/EXi9Cz6+ft+hNeDOOLyP61oBhF/jnLqOd1
VKTUzZIC8XejG4yM7TE2Q618C0GmJuk9ZuPX1kpF5oMEf5vBn9jFZk1XKtAvPriw0cvymfoHDx2E1l22BLE5AmbA9g+6mj9J2MAO+tmUcbP18HUPOj7gwBpN8w8gZ/w5
iziYJpH2wc2hvJfPCqQ3xbrYkugn+hzTDeyjnm37lM/mMYlxpK1H8H8dLqPaifMfJizoGEV7kTm56598u3M1huaCH6xq8a/pluVIuo6C2bwcAd32Z5jqamsaDmebJBkk
rHCVl6PpVRLjSlEChJkV64O5cMhp+JF3w39h0FylH+2cX8nvCuaiz8hB6qJojiFJqaM8hnoVbYD77wbj43QE/4+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cIbGC9X7iR04g9uOrJthVooVSe6Jm5FvdP7bXDjcNMKSY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwM+piWbBB3kYcqyNQWRgtSEslTeeB1qppym8COwKtpyxM70m73oHsV9CXAhNeYsa2CVrOw4WGbop5NZFm9WkaOaopknx4lPSG5t8q+y89fne
Z6uWUjs3FyzWYQgNX3mWyIe46s4mPnSXDNuOR0DP6mc9e+6v32+1u806mbJ+Sz4NKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwHtHX4lEn1ezQZQycNB+ByGB73BKmLrFttOLcyaRjfgsj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
FCgp9v6knUdJR0mjkoCy5VdKcHpIKg3PX57dHrV3hpfhBAOw4gD1gY6OmVOmdBVe/4IyFdmzkshj7nKBpyGwBFbTISv/leywyDT3xBQKrLFAdn70W9MUKB/LK8IhHpJa
g2BYkH1zLVK62pcwcpHRMM+oJpXGO8M1XaFPvv9OfJNzg/aQ40eCqyQaxBGjn3HFj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
10U+WR2lgN3oGnBGJmtWMqh9YvXO9l5me1DPZ/k1Ji7lEcC0J5DFL7H2YVwnn+TOj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
b3goGvMH8ReL0LPr5+36EyB5abW/CTIw0O2H45vrf6UEOE4b+vE7K+oMMV6NZJxHbABptEsVDWj7Sb3o5hOD5g3DtfjPsZGNHxgXfbwlO9T8wBdJgAilYkTEM5SaWdH6
lK5CPudhvJaVhoDl0Pt3IedvuD7i5X5++7BJ1jsjIAcEOE4b+vE7K+oMMV6NZJxHyDysbhx+1hpPQ4+mKfqlUagoGgaeySJdtTu2QE6KjiuEpav0GmlUtsfpXXPh6IM3
lK5CPudhvJaVhoDl0Pt3IdvRTlztiZVPvC7nuf+AUJAEO97cRgZd7lX3e10IRFR40HV6K3htE23hUSM439gYwcjXJZc+cye6nb8Uj4dRS3FQ6se8clDGItyfREQTAn0n
EYs0teQc5y7Tf0jkFHFCrjGqLdUSeobGF+Zk/ukN4Vtvi0oQZT4lOnHmelyddK3A6En3sS633XyD959wcDCOHhokgsYpAC2fg2hvoOeH3xQctvtP0AllRzystN03E7Z1
D5ofTpYqj+10g91VjPdLlUySzzO9r54718P3h2LHFgx5x3EaCYltXHxeOi68acmfLaYKRb32ITljq4To1ZzzMQDUNsol/KLGhQKiT8Mf9UVzg/aQ40eCqyQaxBGjn3HF
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA10U+WR2lgN3oGnBGJmtWMr/yvTesxDaSNXcVVer5PgmuyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAPEr2j95IPA3Jrmu+FY9HFmaI5+U4cBXnuG4NxsK5QaqPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0W17j0ZPQQ8/CmNW71yQhVIekc+J1LmMqhdUj+at6o+btaAIIPQe9ruwHF9aMqTLb
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAtk3pSHEJheRoZSDKh4RZSbKgwvaikSdfcgWrndAcQhOqnUiNVfi5tDjveir4U1Fm
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAvxJAmMIHUzItVBpniSmxfEuRxsGkXGYI9IGJm7bBp5DsPEC1+g3SeGvXyJQsDW7O
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAtwS4EiK9to2zeIBwToyI3+MPCiQGk1LzRpZIv8qm1OCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAvvWIIJanZhqLlJt2oDeHCD3n1nrf/sy1wGOncBObUMyGaiEfOZw5vTrecEnSUc1KuyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA56pG74h1OkOeSrTdNGGL2V27dBxsbgH0oJNeCejzy42im0L3hoDT1AeoJE9b56os
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAJDeIOxrbpUJuLuoFWLC4dyjB45bpHUM4lW9Yc29yYoGPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAXwxMrjMhrcHwVM0Ew7yAJDoW5oIPmDoJARVoHBikjYwm1LtFlptLBuBFxztlWuwoKdmWUl/cATARhimBO1d/L
ZLaNWFCnPTg4U9Iyd/RHz/FVK/jMGlCY8pSm1nYE0k3mcXBaxWZoU8r7fYlKA8Csg6hRqIQWR8u25zXquDvVMBpBW4heQEZ38tugPAvnnRfUbXsijpgGFXnF7jm6Qy1z
/c24H7KXFBB4WokDOIWA395jqiY3eqNFZpxXiSJhp8diG1tzCg9zMGThTn7i7LYAfSPndd4pozGPM72RZb5OsudYUxIpFFmdDWC79w1MTNZBMDANK/Lo+bcp88+yFgRi
cvkeZXh2YVdMBGuqU3WxRYn46avWbWILHY/wUHH0ZWNxgoJ3oRtCtw8bhqgEsHrSBZVaYe/+wf0Rud5NwCcqgzQ2Is8uYpTJr5aU8eVOhWHEJCx+ffwrePZpuJ4beALK
CIHLz4q/G4s4yXgFXtrZ4Y6USP8zyagYUS76SwW9SAV8BPNLrFgOdX28ve/tRP/4dsqeuQbQtxBzfG99CkFYHDCcMI8DRGpjLxblPIosoD4zpa4H89fHdS9blfEVbtAy
8clmvy+o3wva7zUCHoNlLmUIFG12VWR5GFFzK1itYDj7fe1IhpMotDCH8MZKRgcVJhbCmWl2ZStk44jhZpYRUxUH5hM/VIEr0jf1PpdL7yiJ6gUjEoWRxT8O3/Ss/Lg7
W8vopTXJFJ8dNz+c5KT/TuQyx7Mhrlwuz7ZLyxdPP8wEr2T4LeT6i7yBRelEQWQDUfAxWBPrPorqdQdRV6p+RcqIJtEmvYeBjKtfeWMCbYgERNeKynZfa5VI8QAec3N8
ZaHBlVrR7dLACwpHaU2PR8qIJtEmvYeBjKtfeWMCbYgfmw6BiXQEzvTHXJVTxjBDbdhr+6rI27LLuJ/kpCKdd67KornOxBT3V7fwqFO9NM2PtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMDchmw9g61ncLcS5toRa7giZNg9p3dkZq60VmJeVO2so+waSwuOpYMTK5kdbK2xfPOuyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAb3goGvMH8ReL0LPr5+36E7iKjn6HdzNz9hDNycNcDCvrsgb92Z1uMP+pIVsWVR6h
F2ctBvXw8CIdQaTgr5YNGubAMfb3/xV/5e0jOUaEi+WPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
3k94tTdna1I2SO0r35wfKoMiSIw6ZYkC09v/l4n6ygePtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCJE7Q+PiUACXSIrCdNk1uM
e3WUa+BrZ2dncNzN7QV7aK3/wlgnJS74dI3Udpk9F6LofSLYcpVhJqx1ut1YkytMZiq/FL5w83wRTl8M6P91OrR1/pXjQ+sA82pGNwg34uZLWcFToSVXQZLT8r0WGsCE
YU66L8hfB18Wf6cz/gAVzlf5jbjNcb9xwpMlAqJr696JGCkEcdzxskkWxam41yJnj3o1eb1oIT0I5DwMlhaJC9u8ryYrGD7R14PwRoRWH9nWZ+y7Gu0mM0ApB5PT6kV5
YpMoCy8Yl88lzwlON6pk32D9XioV5SMTqmQg3a54kIQ6+HH9/+ulPjGnOF1d8OmDfs4o32pAxjamUknOcrk7HkUovIIEx3iXUEr7D5JUOXVEnCcqZ9OM1wT94wNQYO68
JX2udB13TIyXSRE5VjrzOlzwKRzqmIkex3QfTez7T+s3SQdtSbeXVDJWTq0O24u6jmdo5/pBibwms7hziLsc5eDt/rlzEHw/tu7vvg9GvRcCUlkF3kvqDwi1FZl/KqwT
CknO6q/DAdTNWXPUCEuRwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwHXVeH8r/BWadEgLeJooSmXEM3YNjOwgUkFS7jy7S6+r
4CqGedDI5oTaLtBJKr9uSQpJzuqvwwHUzVlz1AhLkcCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCLCkiIoFQmWqIhtr5T+nsE
GKzyML/nPP4x+5cy6V67N3va5oWbxXyK5VseQbkm4eUZ/KLeegzBACsFDRFPMWmHjSsifLNaeP7cRtD3NJX64DF3pUqK17a983RYKN58LWiJ8/Mf5k5qMp8umjP6QJ4+
q9n0r3AEGZo9ilvbnaWmYTHOZN7CienL9anhhkX0l41LKPYwKRgLunob5k14y5N5eHcDrnW+nACRip5NED/ztAke3ZWWBFsXHPIf+Rf3Hl/KYU8u1ZH57YqlNlPfhyNC
a+Fwbn/iYQcrOI0KYYWdtasKU84f7YgFMa3prU7Ur4Jj9FVjcs/Zenudp/BPh8Tn6Db9PO+COB4xf+nSveuqR/OE3tWxbpCdh4x7MPaVdFK5nLbd6simEivQ8J36MZAH
IlvHTbtS/LmJztw76G+DoID8TMcSw8cu4jrt3iZM2jILNNyRZ6IoEFujKBb+mlteTwZ9Y7GrUufUNjSIxp5dzCjB45bpHUM4lW9Yc29yYoGPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMBL+Lt/MJ5cEBZMY0HIEqVI7oH2Ju18JUh9s0Qzk00Nj1JBrIlVvHa0cjxhz/rbZIvChL/R0gMkCGKpQYDa5cVQ
KMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwHgC8BbS98xeV9WreJJ2PkByfSKQFMzRLAFQqYoGXVJy
ytjt5f/JP+X9M9aVGoup54+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwAHqOIDXDuiPGqGsB0P/Yr7MHLgP9XprzpFaN8dsW16t
TTsbaBG85MIhrflncV2UeWtAKlMSqGaUwJ7e7kWiPYoiiuHhDf9ZMTqwCl/Uxj9rj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
3etXJmqPPQEDC+mjt2yOPz2ebzwCUIuVSEbiaxm5SwbrCcUiIg1qpjKsZqHg3jJASyPxTpU8OYO5qu0ROpCuvI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMDRA9Wgqir1roBWdVxQuFrgfSPndd4pozGPM72RZb5Osi0Rd3nOZGnqv6DQ0ChoW0Qfc7jRfMDvrkR6ByAIyeSn
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAFCgp9v6knUdJR0mjkoCy5b8Na3zBMWsc2mxt6EliZ7F3BhOteAbydgFedXyQRBmh
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAHj7F3Rz6xogmkhI/T6QCNGvA/CMn0bSDT+dr4fhrfhxYitCQ+TUndWZ8AivjojCo
rsqiuc7EFPdXt/CoU700zY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwIsKSIigVCZaoiG2vlP6ewQYrPIwv+c8/jH7lzLpXrs3
+aUhBeCzpNnAzHK4eQXzz66kOpCf5tTsL925t11pbW+uyqK5zsQU91e38KhTvTTNj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
EQ6o7T/L8pIprHauSdd4DSn1wwV44acKYQYbMskzWqSPtagXLq1tG4NLEhvJKIDAFCgp9v6knUdJR0mjkoCy5d7AZY+UHmunf8IKdLNF0a+6oV4pNkolWe3nFCiqQiic
KMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMDzBc0tCsKRFUJDp9JUP3rP7chrW9ESAjoOdTw0suyGOYvH9BXI9w47FB3KaqIVq/sgSYyvVtufLF5ns0ScUSSM
c4P2kONHgqskGsQRo59xxY+1qBcurW0bg0sSG8kogMC74w4wEBAepOCiQ0nq3dzKcEARDUwEm7/5ltO3u7bFMckEQGAgtrNvMUgEDrrXfR2PtagXLq1tG4NLEhvJKIDA
Hj7F3Rz6xogmkhI/T6QCNDF3pUqK17a983RYKN58LWhtLLsqjye/fQMZtepIjqSwuBrf/3sCX2FdCpjvyRfbw8qIJtEmvYeBjKtfeWMCbYgrT+ypgbiTRtg1cusdn1eM
kuJiQaSNrjHt8qz8Vx54aUZHUwVZXNSxMaY+yp20hjSFmo6CiOS9OK+d5UfozPdNAWT420vr4WG/TG5E2773Ibr+NT3rD4QwM7MsCSuyj54ktmkIAuYDzamekb1iNK6U
fW0udwAgxIQUpIBb1Cqmjh2fOmKqpCQi2mYo6ZgJgGCu4jk5gW4Ilu5x+kQnDlz/1d6JlEeD2G6sNbXIQ5zFFZLWvpoUvN7qKI10OUfgSPymaeeOBNpuIf5O9DJyW8CD
wvTmkgt59FHUSL+m31aTz2GL0ViS/C2p2MQ/nlIRTFKz4rt0YjscAQEqVVZzgX0rPn5KXOek4dA6f7ASHCRh65ePJ9P5AkOam38wAj7RGRAxAKPDlXAPoJu88s58JPAm
OYEkBqHKVWvku3j0lhr5NYpPZWLY1b+WbLBAiCmlYGHTAG/2ZiKfoPbV5aepJpDS+Ai0/MrnZzkW+fGBOjIwixALGSDMp1mc4UaOBfTXUG51f4CDwgY0/P42G0y+MEld
EO/XYRKe82e0GrZCiAkDxu/mCcYfV1WqI8Qbo09h56WkRjjzu8tCtBL+Mje2BRsI5VIzr3vauohFU3aZpfhO7IlgLXrPGCyMjwkMshCrm577NzeHP4zk59IGYOtAiAeN
ahuGHWABwh2Hq9auA/2eRccp8UR1ywOtnbZ2c0OxBvcmjP/ugYLEhZyocOQm8XeVEPauEbywznWoN+q+nbTfIpx+7e+P4eF0qz8myC/v7y1yfqyJM0z+YSMOm5UYipI2
LZbR7CMG62DOmoqfCbOaUebkecC9P734tBodsdJjwd678MN05qkTaZfz0k9wP0cxOEGmQDr7FVvpJP3TmFP5XyjB45bpHUM4lW9Yc29yYoGPtagXLq1tG4NLEhvJKIDA
my7CbUIeRFMBgaIwGoRUNl4vXuFtRPfG6zBKoYci8DQ4QaZAOvsVW+kk/dOYU/lfKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCbLsJtQh5EUwGBojAahFQ2
0rIDmDZwbHQV7daIslkiudPQNDU/3oZawaMDNnnOgAbnL6UdBtRtat0THdyTWKMqj7WoFy6tbRuDSxIbySiAwCEcKctpIqpOxoU6RmfkgoMJbsISb5b5flBLArxYo532
t0qTEyf1Rd96xWiLMJ1c6hZNPbXcT8Ss+w5HzhdQPKplqoQJFQeaqpfz//cyVvtq5y+lHQbUbWrdEx3ck1ijKo+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKD
n9o8OB4lxgdZCTgO7hM1wxS5Mm8ROkheh/y8xrnRVICCJ/x3L82rX1LdzZ9kM9Nwj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMC5ZKmE1yfKOaBYFmeeksh8
Fk09tdxPxKz7DkfOF1A8qlcBxNdpqD4Eu3v4fZaThaaLPcsawhLVCxQ5gLueKRDZVU1iwvVsmL2Rgra/oPMDWBxXSkKAzBa0DlYXNlj0rHRo2MXqxCsCZNX8MXsDFsHA
a4uRXgWZfldEKfU6zDpi+bDSX93OAnkJ9p6LW4zFiQBcoLDpXYLXpiSWzcgZQ1SzpdvtK+FC7On+BuykDmT9TxUH2JGveZQbgeXW78T1YQBN39RqTIdRxcUYrjWfkIdK
N2CTQzrM13eNg5Y23/sDq5AvdhUgmNUhcU5ZjaOafGXhueyVNUk8GGr9KFkldZV2fewnC117WgpJOY0EwrELO6OgSRn9X07InqLshyoENZX0a3fQI5aRgzxP8ODkgoEz
DjbpftV1pOyji4sUb5LIMLpigdWkkPlx2p0yP3VbsDVYojP1D2/DHhHjjZNzdsmvWBFludW6HmhSw+zSThl2hZVulMIAT6wdf3lBrw6ygquT9BQjXzWIUtt4lIInRmnI
mCc9TWbOBZjeCJ9VmDvfujeavl4S/YJlbkJkfmv3nl1/NryVeNYPw7qSEYE4ON+Ogif8dy/Nq19S3c2fZDPTcI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
eNfrE/+ntCFv0/81692uq+wJc5eL/qTu1OT16HEpUr625DK4207nQrojviTuW4mPj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAeJC11G0roGmLHH9VqDw6r
7JMGwBR/Mwam5WXlEX/+6xhrrvALXR7PDPDmMtmtaq0oweOW6R1DOJVvWHNvcmKBj7WoFy6tbRuDSxIbySiAwJsuwm1CHkRTAYGiMBqEVDYWTT213E/ErPsOR84XUDyq
SegHBbczjiBHQUHIeGFSJcLKdNSlaW4YgcbBnKDRkT45O+q8jsiGDw1H8T4YXFyiFEbxH3i/XStKpO7Pn5skYN/Ks8GyWl4jcSRqAU9DC/wZYaROEes7FT9ol31GFPkH
Fk09tdxPxKz7DkfOF1A8qiJM1Z6fzeBL9txoQi01WqlMd9GM7Ntm0mIOqATt3orHfNgrzi/S8fEZDhomekoRUo+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0
n9o8OB4lxgdZCTgO7hM1w/4nArHZe+OqzAlHDxmG/kOCJ/x3L82rX1LdzZ9kM9Nwj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMDsUjm/EBdJLc0o/av/3kHx
cTGV9OiO9iztSM65IPWrlVJJW4nKgMXxurHKO95HqW4QtntHvUJlJ8kbIHopBHUPIXQkLYgFVVq4adXr0zhVGLYSdMVCmzQFSGO9r+fd2Zj2nCSyhQmK5+ohskrKRpeW
0/P9Ov1PeMtP5c0Suw4Dr6h7lxwRc5EEFUJ4nFt2nhVZJlBVn3T+aWr4RU9fq/6xadWdk67DEuSWDO5p94k9RcBAcLj065rF5slmRaGbt2ttqzPb2WMSFIjfwjHJZqNE
ECKAXIfeTf8T9iKDwA4eO4vv+0sdQ9IRSSIe0MBUl3uQsuoNBMFG2d3S+MfcyTVOiWAtes8YLIyPCQyyEKubniyJWpjpgNtWpCPV7hSNdSs8aNn0aBCHg0mjdFO0QyJD
miI9362LMLPNZZ9m2lLDRmJu4OJ43r/pgsYnaHd3zJIKgpLgY9H/RmbYcu0ZfGWRqSZ3kT9vKMpirinOSr3oFKVGfhTeil6Fe0BI3TIUj8CaIj3frYsws81ln2baUsNG
0U9fALl4aZET43e+xLTiQXOD9pDjR4KrJBrEEaOfccWPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCx2sSmoPfMrQbJYSg92U0X
oROs7QItIuZjT+zPkd1aso+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAMd/E/WoV/nLDWGFFGFqbO
OWk0W7U4nobfgHfGFsQkw6t3/c/QRvKo+hLDU0cOOg1zg/aQ40eCqyQaxBGjn3HFj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
yDwLQG/E3sfimF0Zm1rhupQeufs+guwDu0syo9VqgKmIEOiXK2dTPlsLOA6r8YpEj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
L71iCCWp2Yai5SbdqA3hwnrwavuw2YSJPhFgU++QdO1jwohUgEohUgoxpZTd0Vmn0L20LJ6GEl9WYyR3RAp7MI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwN3rVyZqjz0BAwvpo7dsjj8l7w+BDeFpJJUEFA8G0cPGL/bouRDBLyS/qzQftHNXL4+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwB4+xd0c+saIJpISP0+kAjRkHfFLTQ6Bc14v4r+fm4eicAPEOE6Qn21qbNBlTaRu73OD9pDjR4KrJBrEEaOfccWPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMDIPAtAb8Tex+KYXRmbWuG6EYkGhoSdhnmNURf99Q69J6qdSI1V+Lm0OO96KvhTUWaPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCesVbDrkHQ2Q2O8V4KCnvA+p+sYo4HI1lhwmTQZFbZnCHjHq9okfITs4dkZHCyQdOPOxsoSXj+yWk0yvwujJ5T
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAGeaCSKLJtqBzjaG27/0ZBE+w5QjoOrBFzwjKa0tqg8IlaN1rmPRd1MXqNMf+wO52
EnvYHBpSVf9d9lPxQ4kC0Y24fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMC2TelIcQmF5GhlIMqHhFlJ
HWQZFzLnJbz1vO/p8cMiZRumS1NT6zsbM3ABpzhK+i08+hw+O9OExi3XPO516NcRc4P2kONHgqskGsQRo59xxY+1qBcurW0bg0sSG8kogMC74w4wEBAepOCiQ0nq3dzK
kDHrR0W3a1Uv9Grv343cRIDa4Jtg23omczHULFjsXguPtagXLq1tG4NLEhvJKIDAHj7F3Rz6xogmkhI/T6QCNDF3pUqK17a983RYKN58LWi2aO/RYvR9vbcKqvBKIG0H
DE142YOBuQPa4PxSxCRH7CKeGmsTvKqeOzBtuTlAQXT3WRaT2hAz0gYxW+l+5m+c+B1bsvHZB2tr73zhbcMCkvlCK2Dvux/4vZ24L0hx5123vTaBQMsJ7Uy0Cp8hvgvb
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMABFg5NyA1mlyMaKOYJCivAKkaN+OEwxvPh2e5XbQ355424fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDA
Wf5s0PuxtgTUL8+pRYJYzpGegHjSJyDBoRRvRUsXLUxKoChkJjHoykAbG5R9oxL1j7WoFy6tbRuDSxIbySiAwGfo/hT16ytNQCQ3H6BnXYfpJDvTNs7QfS3MmxYCwZCe
dqeNVWRwrRNw+V4rO29W1KIlRbaQs2Gxx70NHUQhdhAL9vq0FW3+Z9Zzc+3UAoALBSS40ejRl5DYUTbbETxLR8OyOC4ITnSfN7Xf1qyd3gqSBL/ODt4k6IqfGWDnvfG/
hFYEBnPi5Zgz8cxt6gMTPp5hit0Q0l6OIzjRZ0ilX3xiYKWQfj4bbTeeIgMqIrtkzUDNH+DuDYKm6Go1YmkkgBjUZeGnjOquZr2QDtixhb5tIEhf7p1rDhg4BSu2evg1
oC+E5Dsy0uOcDbYup13CnugV9JAd/+Jxn/qeD9EnOWwjZkZKIVfUtRgxkKROJSCnDyQYLnEg5zoWl5V/XQmvIeKgWkFfdi+Z9N0zNilC96AgAOX0PIzP0FnMj5BqYZgV
ZGURaPu5ci3WpRDJknxWu0ZHUwVZXNSxMaY+yp20hjTfrMmpcQ3uAacoao48Wci1sUjY+lC4+H5w4xKUZh0cmjCVERYfknGMiXui5ELloco7fuVAeaSYKT5W89/nVq/5
Zn2Q7srVwq0PBnosfMIkAU5nqFvxVtj4Zc0Kh6y9FwLvxd738U3vV1/EEh8v6F2P5T/RVMnO9u3gkLroBJ/X/cM2tE/rioWNAYDnIA8x6YloNvS/Oz4w69Lb0F6Krd0y
+ckhDxrCO7of9ok7QilEwsBHj7B9MIth8UcgW3vLTOFbGhXGINzfUvGWs/DYIhlfsYy5IRqJqpyUt85u4dpq/0A7IK33t0kiGm5OW+ZAOPSyADDg9tZCpFZXRloCQN1D
5T/RVMnO9u3gkLroBJ/X/cqIJtEmvYeBjKtfeWMCbYiUdBjvN2BrQDR13eNHhs3CkiQ0jkRySzg3NFPTxcsF55HvJv/u8GMKh8p3G41ofBVJld1HA3ixoQP+zzXD+t1M
jjBQ75PEGCAZy4xAQPPuZ3fcFXmxHmpAiFDisW4lBZ4ryaL7nz06nQjyLdLwOV0rhzIK9XXbZZygPyNAlseOfgF1dL6+1X5Ynf48nRE00OjhpoJFDStBKIiH1rcA1r+O
Tx50enQIFzxtRvl3ziPlc4nRjj0cZr8bXY+RJLVdK3PrhWINw9s+9/bVMkhCdiNgOEGmQDr7FVvpJP3TmFP5X1rChXksy+4Op4r7P5LWAsG7XSDyJXZhtF8Dqs34bKfU
sbjbmX6R+sr13HgcrtDcoZK3BXDf15JGYcRCKd0WgKmv/p3pZrXP7IQH0q/mwBiPa7qUG2wYWztP5gDFi5jD/MVCfsYPz/MWT2ZCEWswUlWOMFDvk8QYIBnLjEBA8+5n
kZ+uAFdzZiEr4L+ujCLSroEt5P1f1yAaIBdyBX8mC+Hi5cm66f7tBitPxtYKUakfbaU94F6UqH9IkDi+cYFrVhlhpE4R6zsVP2iXfUYU+QdLIMmzN/OdAcTUf55SO+zt
tm/Lzmm5I26Jt8HuvRTL/5L7B3skzyV6V0aQohkOYQSBVwvbDt6Fr053WLHZ/Hsyjf9T5tRnamI0Tmz/Opc7EJP3BDlr/nvSTeyT8s5WgoG7yogS0VCTMEXfP3sdZDG8
QxvdQoWsLxJu9tsNWFXml0bmmiT18cnFtiXxCvkyKu83YJNDOszXd42Dljbf+wOrkC92FSCY1SFxTlmNo5p8ZRMPsK9bMMbmg8qX2ui2VzzKiCbRJr2HgYyrX3ljAm2I
0K0qjM/iqG21cf1aLXW+KBgTmLPGbqqh2V77YN0pyCvg63vBxtKqQbXhO+GyVYSWyogm0Sa9h4GMq195YwJtiDhBpkA6+xVb6ST905hT+V9awoV5LMvuDqeK+z+S1gLB
u10g8iV2YbRfA6rN+Gyn1PVUNlUNjX/qePR8gsM3+RbsDU1YGNBFjojAE+DxX04/mOJ2N3017BJJZr1YD5RSq2kBf1Evh72MzG0jGcqym9nV3omUR4PYbqw1tchDnMUV
S2EiOwH5YMNzkkJUIipFIxheulNDyJutVqJ8aat3mDcTIWCRCrT7D5wBkuf7ew5CYm7g4njev+mCxidod3fMkgqCkuBj0f9GZthy7Rl8ZZGXMHbeWm1IG5pxdn1wntsw
q5WIqvsDhxh1ODDKupRtrjxJ1P/ciW+fZJQ5ZZbwQASNuHybzCCVjbv0GSSWZ4QAj7WoFy6tbRuDSxIbySiAwOCABLjGX+83ZJjUdyx0FNvbLBOP9Pzd1AG6qUEjyql3
7PSJD67dlHkxZ5qJ70R+P3OD9pDjR4KrJBrEEaOfccWPtagXLq1tG4NLEhvJKIDAHEOiJYubEiX7CvnDXKDZ3G3PlZqU0bgbSOknSEROFapPP8UwYcRqcT1p0FVmUxhT
qVude4YVRSa1XUY8wT80QLQH+8eTWiWtxV5Fqv1apXhXmRClgRcJzrOkUEwGlMeo39rE9TIn1XxgAeYntGrxUZkIhsjiSI5veua+gwAD9YsDWB1sI35cg2VA+xtpsVn6
YdoHO3hryDLfVbG+6EzPQWvMZCXfj4njZjG69QGrzR8slvYX3ApOCrRaeQ18lITPi+/7Sx1D0hFJIh7QwFSXe3wzulXowbwLeNMmJJkwBQkW67/EFqTQLwrBDC5ujCHZ
sRsSUQiPLVWFlzz5r3lUmnD8DRGyAcMKKx1LnAozYiH76jB0XKTasgRWOT9xOXA10XqG3muFeVlsIvK5fycYsa19hhBemox3sQDbF6DQjEg0K+yo1olyeZNhtpcCFHyP
jjBQ75PEGCAZy4xAQPPuZws4FUTQ08rlNdyROK7cWK7RlgZ6He8fHkV3jn4r6L1zFcV2x2jP3h4eQf9uQll5RxXFdsdoz94eHkH/bkJZeUdy+s6b4Ka9Jl6Mrste+tIt
RjF8XJCL2h+ya/t/bOWQ+Ru9WSM5Eljm1t6MHHxAATT76jB0XKTasgRWOT9xOXA1iYSVv8e4cn2QMDOmaQPOk1/wZTi5ihElo8f2QufRYzWGzoSJmD2GKobBToIFUwJV
sP3LbXkaFGQzU/07gT/Rh2rkMDT9kUW9m9lye4DzVJ+lxXUO7GzF8xDNShenie1j46/o+brHyzTlelK6tf48gFcQrjKoIilvjhKDdDWGMmmPtagXLq1tG4NLEhvJKIDA
9p5uZi3Tl3upZo4/iJCBl8OWmRErofcUpTlaxMon2MZm11TjRVgCBvAXOxUjeWYRj7WoFy6tbRuDSxIbySiAwLKDsr4oKygtbg6zqZ+nBsCcfu3vj+HhdKs/Jsgv7+8t
l2huKOpkeRtj9SOXia9RyfvqMHRcpNqyBFY5P3E5cDWJhJW/x7hyfZAwM6ZpA86TSQu7wxTsuUmkMGt9B1cLk3SQC5vfaCZW1iFACuwqc5g48ElFOZCcsHuLMpZoMpWR
1YX4FkJpeQhDzmAsmqZGR4lgLXrPGCyMjwkMshCrm576Psl3e3m0NRtur1Ag0HyTk/7kk28LO2wyXU2hfFEITYbiGdIX/yzIvYc0ZF7BzufQUIkpedahQeByoXe+DLAy
8b0qqSjGDgcV77iDxmUsdHzYK84v0vHxGQ4aJnpKEVKPtagXLq1tG4NLEhvJKIDA8gbpHCSRxX5UwRhegUdhEQC1zbHJnMJEtNH4S0LP/T9HkjyvxNATgX0MMp9qRGZj
CknO6q/DAdTNWXPUCEuRwIkTtD4+JQAJdIisJ02TW4x8NO8FWCfdPy99weuUlyT9JjdNb/U5+KyLA9OAZU1ZBiD3gJnAkCeAlSfiQ3URSo4DcdmOeyAUtPvsr1kYw1bl
arWomxjfodCBOPDsob6Zf9eno+JPLGypyrnw6HT34SSt/T7/g1yjC75Q2dWng6t+bEfWCtR5jS57zqzg4wM9/+UBEUA5ixL4ZpunzF4T25yT1M2ibCj5CcbTsZhc+4Uf
nTd/m1ZciEvglsQuUNrP5/aeWiwJqug1kbrDmEyVU7tpJtpDgHDtebTFiMKTFmGrX4mHlkoCpt32Qqjew2pUXsqIJtEmvYeBjKtfeWMCbYjIs5ld2fVuZQJJdnzgDkvX
JQHrOpH7paML4a4BtObhm5x+7e+P4eF0qz8myC/v7y1r9ij9YH5iDxDwclztZp8XIzHl8K8FJvRHhnmVPaD06/etSo46JNIh2FMgyDkdWK7ynTFmY3pQ1PkTuuPeJCIS
qHRTqzLfmH6ZZb7Nyslc7Y+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwIkTtD4+JQAJdIisJ02TW4wBnziDHcuPldEe8MD/0Zqz
9OsUJlK+kP7GJzlzXSSsfa7E+9X/c0w1O7KNEB1RcfGPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0
OOHJ5sQkGp4c2k9q6VYiWg3dNmEcGypOkq9KocD4TpM1izt/kW0znk2JZ4FyxKbs74nlmR/4QZhe/WSqI7h4fI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cLtaAhI1cBHpifz3NLM9ExvKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMAmHbIsy7j2vbBolihoIMRX
qbS6eW80NNMzwfQPCtZxxucvpR0G1G1q3RMd3JNYoyqPtagXLq1tG4NLEhvJKIDAIRwpy2kiqk7GhTpGZ+SCgxAZrhHukDjY/Vs1R0frGF3YXKpuZuCG+ysv8DN1fdjr
V18TW7qmE393fpCUXJB1lT2+jGsLkTP0eynfMABVY1fwt7v5LHBpZo1Z9UKNVycVzicFzDHaZ9IOVrCE2DsBImFxUUIJ9MO6FfsItJ+7LRArKo+rTSwJtr9ma1q0KlSJ
i8f0Fcj3DjsUHcpqohWr+2QkNLU50KRcmjfW8Xg8Vi1BmMJYPP7FY2D9tkD0ExHVsmkmal+ty9GUEUpX+BOohY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
DiXjSWWTT736DgBrQfHCVttbq82/O0amnMHdVGRkbjVXEK4yqCIpb44Sg3Q1hjJpj7WoFy6tbRuDSxIbySiAwMzOJ13HROhAr2M7jFs4lSHngk47Cplfv78LkUVK2+zq
2OssAmcGAU5DfkQQs19ZiliiM/UPb8MeEeONk3N2ya+mO72lbwmMEosaVo6EyFYoHH5viUjps5g6OveUhhgjBY8DlpafHZJUdSYDJcsWqI5prmcJRd1zLQ9Z4UG+woGn
WzXU3PazDsKyEoFITyPF6tGPyEFvZ5Ey/g3m1qD1R5SmtE3JZUNFbiGgLi2VpAgY7WCQOVEMFRDDSYGavBYJz4sYEeZjdkPVFsSbzTPhBrv/ALDxn0rDA2liWlB5d7+/
BWsYpleyjclbwUrkJJzjnu1gkDlRDBUQw0mBmrwWCc/QW/PsgpgAgA1zvGxOE0aSnRu+6k9KS/9uQT10PQ6gcoFql46K1oLpPGvkm9arxb9siPdwSGh1oj6qJCdQQkbX
FFC9RJzwd3GF6Qg54Hf17KHZh1ygc+30pCZENmzWlUyHCxksaauKO1g7WrsD3kh4EsmxwXdAXlL1NzWBPodYXIiuscEEAGbGt/7u4+Hxttw3EDGiCLj9ZFT0AIX0IQ9h
f+1vdbuHnskHcZIA4zou0whW+kMAkvF4iw6wYTpcJeO0A7crohYhW4Rtci936VfUYdoHO3hryDLfVbG+6EzPQWBbjgOATkgY/kxTVZSOXQUN+OhrmRSggNerlUy0BgRt
A94Zyqf9REzG3RXdUDRDR6o4rOcRvpiX1bQjMCYkGg2OMFDvk8QYIBnLjEBA8+5nYqtMmuOKAZl/xk6DrOmNGb5xpVV2PRGZHsDnGntBhlOFE4Y2xc+s0SJ3OZuoz03+
eFFYEHOuZi7L6a/u3vPGzSrw4aqLv8rezIjtR4FLu4dq5DA0/ZFFvZvZcnuA81SfrFRo4hSm1L/GHp4mdHABgViAKS8JotSRhVXlYrB6ZtoBe93VtLTc4Jxt7YK9qdrX
ffFL5AihhaxgUVvxl3gQGecvpR0G1G1q3RMd3JNYoyqPtagXLq1tG4NLEhvJKIDAIRwpy2kiqk7GhTpGZ+SCg6BoxC7YXqu7ty0qCrSTcfKXBkxFeaE6HHdraLzf1pZ/
jjBQ75PEGCAZy4xAQPPuZwpJzuqvwwHUzVlz1AhLkcCPtagXLq1tG4NLEhvJKIDAd0BJvQfSoQx63oWdPsxQQBFudugx73qzOUOLqLO5VnS6T2UuRsM/NoYSVhU6Y+18
dlN5ockGbu4hC5c/LGj8zo4wUO+TxBggGcuMQEDz7mdMQFFHQMJh+SjaDH6ffJYdBP0eVwTaI/TsSRbzgu7RWtClqBYytD8gwSQWU0DD5zEJbsISb5b5flBLArxYo532
t+F5/xx6nup5As5wWRkYLxZNPbXcT8Ss+w5HzhdQPKqBrU8GklwFvINYl9WtA/875y+lHQbUbWrdEx3ck1ijKo+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKD
n9o8OB4lxgdZCTgO7hM1w/4nArHZe+OqzAlHDxmG/kM4QaZAOvsVW+kk/dOYU/lfKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCbLsJtQh5EUwGBojAahFQ2
6CT7wxq97a/RNBJrPH4FgFCEWMLsJDFy9YpcV5g4+giZr+xoG9n7FJ47BbqqrcEZOYEkBqHKVWvku3j0lhr5NVD5fjvdTWEaKUpyu3j7rPB9XbXbjyjkQvbhZGIABTsO
++owdFyk2rIEVjk/cTlwNdF6ht5rhXlZbCLyuX8nGLEvcv6u7V2lFfpcEhQKGTaNCUcdQWpZXcaNeSC8R6xBsa0Xt71K6Gro+H2n7fYJS7L8CvFL9nXrqXZvAioIb0/7
lkI6yO1Vbpz4zMNAkyr6cFDjvOorKGPjKKJi+cEal6/BrGRN3IlqZnD5SsZm7tPkcCLMU4paoJxAK0vZJ0DnmxlaOfbn/fARKh7r9KYIzDGPtagXLq1tG4NLEhvJKIDA
iRO0Pj4lAAl0iKwnTZNbjDhBpkA6+xVb6ST905hT+V9aJGaCZJ9xH7s+vZQPfiSZ7IFCsA9len9Mue5bNVx1Ne/M6fhy60rdTssODU26soCuyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwN93dNjrBrnDvi14iMtzHblAANe8w+twOMbMmUQAb5/TM6doiVBguibNVuoafYYbhMXRQt6FIGCbZVvnxGLNj4RprmcJRd1zLQ9Z4UG+woGn
++owdFyk2rIEVjk/cTlwNf8SlWba3mkMf7Qppcwuil3+DRvIZi/BAcuJhkm8rDZE8SZtwoHnq7h+AV6QJDMoKAPeGcqn/URMxt0V3VA0Q0eqOKznEb6Yl9W0IzAmJBoN
jjBQ75PEGCAZy4xAQPPuZxRFMGQjhEwyZYuZPgvSC2boOyeXxGJzCyHRXGsR7htk8TMJwksAznUewo5SS0shI3l10lul0hi5Ot/oa+hAOHJLx8wW5qZRicXuMYYeLqiR
wEBwuPTrmsXmyWZFoZu3a8qIJtEmvYeBjKtfeWMCbYia/7eDlVPPvUBtZxxfnDwuyogm0Sa9h4GMq195YwJtiJx+7e+P4eF0qz8myC/v7y27MotcZIrVnkJpr16yduMr
ZrWgMXTTNFLghWYRtRB4TY4wUO+TxBggGcuMQEDz7mdibuDieN6/6YLGJ2h3d8ySzgzpjnEtgIFiKbWYCjxWZI4wUO+TxBggGcuMQEDz7mdbNdTc9rMOwrISgUhPI8Xq
yogm0Sa9h4GMq195YwJtiElmECuKBYJjKmI03jjRJ5TKiCbRJr2HgYyrX3ljAm2I961Kjjok0iHYUyDIOR1YrgPeGcqn/URMxt0V3VA0Q0fJf9tscFxs2Gvgd35plTY7
jjBQ75PEGCAZy4xAQPPuZxXFdsdoz94eHkH/bkJZeUdibuDieN6/6YLGJ2h3d8ySL9nRvfF7f/br0BlPTtS2T3G1KOqtlrcsGnPbee3q15hCZQ0YAvmDRmDi24ndKyot
nH7t74/h4XSrPybIL+/vLbOOj63pXDwkmnP/jlMGL/CKOccL3mo7yWJxEODUP8HNfbNwdpAUFQdDm/cb9VZdMEZ7J0wx58eMNjT6i9FqMcDKiCbRJr2HgYyrX3ljAm2I
WKIz9Q9vwx4R442Tc3bJr7gBk6kxE1h6YA5r0ogbLZ6MynEfNy8LehzbR7mIge05yogm0Sa9h4GMq195YwJtiGQkNLU50KRcmjfW8Xg8Vi13nH7p23vMfO3HZIJ0kUt3
8YdEWwFsJVsUToGbqB7gP8qTVk2B3as7fpja/iGT6e/KiCbRJr2HgYyrX3ljAm2IYqtMmuOKAZl/xk6DrOmNGfOKgXnvsOOIO0lzwWAbqIsSybHBd0BeUvU3NYE+h1hc
yogm0Sa9h4GMq195YwJtiGi9HhWDOuiKNQ0rfwD0NjXKiCbRJr2HgYyrX3ljAm2IMXelSorXtr3zdFgo3nwtaMqIJtEmvYeBjKtfeWMCbYijii9B9Ib5BEfYA+CvOC0q
sIUPDlBoVkjr7I4a4bb2+MqIJtEmvYeBjKtfeWMCbYgHjTOkXDuB37oYegkIi+GKH2dpq5BBRIZnc3oO/x2EfZoiPd+tizCzzWWfZtpSw0bxMwnCSwDOdR7CjlJLSyEj
JqEjyaQSnbH47JQ9W/F+8ebxer55WoY0JpEvL4ySUZOpW517hhVFJrVdRjzBPzRAyogm0Sa9h4GMq195YwJtiOeNjqTlC5FqDQIdRP29W4ygDxM5pUHWFgVpYaJN53K6
hO4g/DrB4t7x0Sp5O9Yxgv3btIyFTMACOuD1ivjttnTKiCbRJr2HgYyrX3ljAm2IFcV2x2jP3h4eQf9uQll5R+1gkDlRDBUQw0mBmrwWCc/QW/PsgpgAgA1zvGxOE0aS
yogm0Sa9h4GMq195YwJtiBThOEQKZ9IXJ7ZAGgEcrbEBxO8XyDCigwqYoCu/mbTwAcTvF8gwooMKmKArv5m08FSCcYD7SGZgXWsaPxsXY3cK8SmGy7U3p1eBgEys22/U
j7WoFy6tbRuDSxIbySiAwIkTtD4+JQAJdIisJ02TW4w4QaZAOvsVW+kk/dOYU/lfSsqXwQFWsn0BslvZ6u9Dmo9TcD2xB4HysCZnQvlEZv6uyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwP/sM8bEFXjmHJRxfAPLCYwhdCQtiAVVWrhp1evTOFUYpKR7ihzh+IOiUwjPj4t0VqqgDUxq6UfENQDvVfNrMd5x1Eud48tj0y4RPx8ae8Uw
rsqiuc7EFPdXt/CoU700zY+1qBcurW0bg0sSG8kogMD/7DPGxBV45hyUcXwDywmMCQ5WGNHqo1lSvGCoMlFdBQwSHqJZ7rmEDhsjZ3ZOYRGLaOM8X1v0X/Jj7IZmc/2v
j7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cJVTWLC9WyYvZGCtr+g8wNYkFnhO4/C6edg64vgh+5peWjYxerEKwJk1fwxewMWwcA/2DNe49Do2Efd4n3LWUnl
sNJf3c4CeQn2notbjMWJAOfZWZnrJuAebJKrJlRrJKJJoBp/OteVD88n836aNTPvxCBeBpoHUjFGZIflFUEOBTzytJnIBbfT+pbojE4ZMJOmeMhrO3cPvsj//q0/7jDo
KJtUS/UhV7rB4Y3eses8IxlOBpE5Hjrk+SXMlw6AoGwxd6VKite2vfN0WCjefC1oPTCoJalNaZ1xrldXxGVJa5LrxRojBKiYDIjwK199CluEQqfTGMKNFyQT3KU6gJlw
WzXU3PazDsKyEoFITyPF6saXaZc6vpY/QgZRFdUOPG9tz5WalNG4G0jpJ0hEThWqTz/FMGHEanE9adBVZlMYU8qIJtEmvYeBjKtfeWMCbYhc87IOTcgLSaToZt+lYHjU
JkWMyQjAL+icFCcRSl7/QiibxXJicY8F/uaWQdgpEg+JKrono00vuQLv0b9UaxbSnRu+6k9KS/9uQT10PQ6gcvloDtv8TpFAv6ExypY4sBumO72lbwmMEosaVo6EyFYo
HH5viUjps5g6OveUhhgjBdPdVtqziT2fp3keEXBGQfRshBBe8k/+GKPZ5FZbR3JKwEBwuPTrmsXmyWZFoZu3a8qIJtEmvYeBjKtfeWMCbYjxJ89kD4bjuwkwrWGQa9jF
HRFOGPRAI21hj6GnXyuUWFWWuWh2ydkMh68jr5agp5hhefi9ipsMm2X0ITB+sGtvyogm0Sa9h4GMq195YwJtiGKrTJrjigGZf8ZOg6zpjRnzioF577DjiDtJc8FgG6iL
L8VbIao/0XHwsqD6xNGU1pKWVBvXXiQpKNKX1np3d+XxMwnCSwDOdR7CjlJLSyEjHg2jezcXCdumbAjBXj1TvS1u2u3hDKAhDeot1WAo48npqXcHCp3R0MsDfjJdkzwu
78zp+HLrSt1Oyw4NTbqygFiiM/UPb8MeEeONk3N2ya9OniKhLILYAbeWJ85qX00i2RQxtuc1Me5QZjQ+R4cEAfT1S1UrCQftofg8SVPQuDEdYxd/UNEQRGR/E1Mt8OyA
nmFo83c8IazQxWNbcd6dvNv2yrZbIQCHY3y8nboRbUZgW44DgE5IGP5MU1WUjl0FDfjoa5kUoIDXq5VMtAYEbfiMWu7zEKNgB9rH6g+1l+EVT5/2zh000ue9lY5Ji1qQ
r+atvIiwnaZZM2cTbYs22WJu4OJ43r/pgsYnaHd3zJJBve82k+Lqqd3+CD7kXuv+yogm0Sa9h4GMq195YwJtiFzzsg5NyAtJpOhm36VgeNStop38LoSCl5t2YrAlofyP
umKB1aSQ+XHanTI/dVuwNcBAcLj065rF5slmRaGbt2vKiCbRJr2HgYyrX3ljAm2IXOa80iXhAn3WlfGa//iTXQ1akmiQuCjznnvj1+DiE55bGXUALXTyia5idSbav9fv
MBc8L9jxTKLCoZD60tFVnIEeoKi4ss+MhHm6tZcbtASL7/tLHUPSEUkiHtDAVJd7NbMjaS3qxII57qv+SYaV2ROfTKv0qf7p8XfG/mY1CPV0eFZqUbbTXIeYIGDppRd2
Ym7g4njev+mCxidod3fMkqjzd71yaZi2kgKxYVqi/9gajW1OSBk/CZW6tk+o8AhUhxDDhfSq0OrE8JiND7dErWJu4OJ43r/pgsYnaHd3zJKDwEKdYuYwF2IQPeupWEgp
Q+tbNLT4L/DNt8ZWdOrzmPXIShOK9lWV8x380Kdk0aExd6VKite2vfN0WCjefC1ouXvH2rtP7KEQ1z/DYFny3/2zM1IzQvw0c18CRMM1hXvr6LEEpd9/DMgr75DYhs1z
j7FaCBm0WI2CGkWqdS1PkY4wUO+TxBggGcuMQEDz7mdc87IOTcgLSaToZt+lYHjUlU1B9FJGQdEp+/s3wIIdEG3ywNRHAfx8IW6ne9Qy3s/tYJA5UQwVEMNJgZq8FgnP
ixgR5mN2Q9UWxJvNM+EGu/YOXjc2w1gU6tZCQaytV0qKayykNAYT5yvrj4kxFQ3aszcrMCBYqjlARpz9g1c1apx+7e+P4eF0qz8myC/v7y1T0/qJGlhaUAwaPPnvckBU
TylXguHHHcU2h2MFSVn3VYlgLXrPGCyMjwkMshCrm57KiCbRJr2HgYyrX3ljAm2Io4ovQfSG+QRH2APgrzgtKrCFDw5QaFZI6+yOGuG29vjKiCbRJr2HgYyrX3ljAm2I
nyY2xvm1aS6sITK/ZUTWfI4wUO+TxBggGcuMQEDz7mcVxXbHaM/eHh5B/25CWXlH/IabIVRMiLf8H/HLuzlx/0MXpQqAUYMWn9ZN+Im1fXP/ALDxn0rDA2liWlB5d7+/
YUXdBK4bG+4oUysB4O0494vH9BXI9w47FB3KaqIVq/tibuDieN6/6YLGJ2h3d8ySbRJhH8GSN1DOAUhQGJLVcIuwFVqZHIxVfToGR35rhZWPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAvvWIIJanZhqLlJt2oDeHClYKclp0BdyDJyzI+mBKzqJWlp59enhiSgwEl4i/cr9SPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0OOHJ5sQkGp4c2k9q6VYiWg3dNmEcGypOkq9KocD4TpPHa398tSSjAhEaJJTjYNmz
ksoo4Df69njFPrcCK/DxoI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwJUqVCNYvATBgTHam5A6It+NHKZcU/sIHLJjMNQzOmt7
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAOJeNJZZNPvfoOAGtB8cJWNnclnn3l6bYqtSQLxxce5lcQrjKoIilvjhKDdDWGMmmPtagXLq1tG4NLEhvJKIDA
zM4nXcdE6ECvYzuMWziVIfQNyW8XUc9+hxR2TZU+pp8ULw5oGejbO3L+EDtdMDTBBlUZi5zrl0oMeDE2bfLDjBVufbPlluZXmNkcWslFlCY1wk4O2BPWGMID5lkEYCBp
QxelCoBRgxaf1k34ibV9cxRFxbHU2DDF3J1Vsblaic1m2riyWpJves/Qom6GPOb/j7WoFy6tbRuDSxIbySiAwLKDsr4oKygtbg6zqZ+nBsBwr0TbT5MEpaBcsse8M/og
UAqIm7oDUSTG4bPXJXdwZI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAnley/lFqKqRcuafeEUotonIWmQcZysYo7d7EoM+XG1MfbFgDAzDnWhWzE0Ob+Evm
YfJffD1YNMST4aW+FKT9woPeyGN1KVB5LsKJ+03VL+NfrEp1LlsQLF5VO+M8GidEsgj9chMYitgYiIwy99AkxHwoeivi3hlRVTx7hiXcyg1H6ZQ4B+aSCZ6mhsrUA/r5
Ym7g4njev+mCxidod3fMkgqCkuBj0f9GZthy7Rl8ZZEUUL1EnPB3cYXpCDngd/XsWj3NJr99bl59jFQzIbUyLQeCdWQNlBUR70y61FsXEalJ2p0TjXQyThndtFV7sy9F
++owdFyk2rIEVjk/cTlwNYYM40zBFKhvpQlaAVvnSYwarkIAj3P43uLs19CVoX4WLR/NZD9PNadsTXrsg4uu4g1YZzbwA/Un4coNhAdkUfcTOTzUQArf/GEc3V+iVLd2
c6ByzjjWDGaV0LZ80CO95/8AsPGfSsMDaWJaUHl3v78FaximV7KNyVvBSuQknOOewEBwuPTrmsXmyWZFoZu3a4oNFtpp0sNh9RPcDppfykt4xptODlmueFfOkMuFYGo4
dHhWalG201yHmCBg6aUXdtsI3AplB/ppvQTZ/WN2KdDPdfQuhXdGn9/7IBDfifuKr/e4Doi31e4BH0cTZs97E4+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwCQ3iDsa26VCbi7qBViwuHcp2S+TZlu2LPv5C+sWLRMkQ7W6nagqCbeGw9KFVzU95+1oAgg9B72u7AcX1oypMtuPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMASKEdO7IHonYd9fV5z2Fx3I+UN/p/VWmjheJ1VvoJagw7hOhUE0r3LKHGJdhdxOadL9hqn8TVYehQuRRP7272T
ytjt5f/JP+X9M9aVGoup54+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwLBcTAe2avwYXw88Hw6wT4fSE9XGF6P7t36TX1eCNg5Y
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAROwsKtxDp822Vhs5FBQuTFN3cC1gD1PdMKun3gXpHKnOD9pDjR4KrJBrEEaOfccWPtagXLq1tG4NLEhvJKIDA
Z+j+FPXrK01AJDcfoGddh2PZFwO0JwIqji6RysXBu0WEpgS2lfPFteXUz5YzOLfTr/yzV07j0mAyMPRvrz7JXy2SQkTqRAPEcCG2fmDsNLWPtagXLq1tG4NLEhvJKIDA
FCgp9v6knUdJR0mjkoCy5d7AZY+UHmunf8IKdLNF0a+YdnaUI931hBCSnDrDotdfKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCUODv/urWQmareFRly3jfx
KUDMxXSbOq0YnhkwhAg2tgf/6wIP6ZpnKXc5CToux/Jm2riyWpJves/Qom6GPOb/j7WoFy6tbRuDSxIbySiAwHhunupN7vLvEaRZOLQP1ZwRHb/NlhhBO3buE1HEkZ9L
m9VUBpci+BeCcfjjQ8IT8ci4f/8tA44wBXJbKmpN3ksxd6VKite2vfN0WCjefC1oBY8ftKyNJRGcuLPJa+avHvEmbcKB56u4fgFekCQzKCjynTFmY3pQ1PkTuuPeJCIS
qHRTqzLfmH6ZZb7Nyslc7Y+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwIkTtD4+JQAJdIisJ02TW4xJVM4qOfPi4u6+6oVGlvq4
9OsUJlK+kP7GJzlzXSSsfa7E+9X/c0w1O7KNEB1RcfGPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0
OOHJ5sQkGp4c2k9q6VYiWg3dNmEcGypOkq9KocD4TpNc0RrTYzhdhevT6jDRg8jc74nlmR/4QZhe/WSqI7h4fI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cLtaAhI1cBHpifz3NLM9ExvKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMAmHbIsy7j2vbBolihoIMRX
qbS6eW80NNMzwfQPCtZxxucvpR0G1G1q3RMd3JNYoyqPtagXLq1tG4NLEhvJKIDAIRwpy2kiqk7GhTpGZ+SCgxAZrhHukDjY/Vs1R0frGF191fJ4lpH0UVtKu/vErgi/
w7Dxs6V8teRRg84vn09isXf14mfxSGHtY0NR+btmCvPnL6UdBtRtat0THdyTWKMqj7WoFy6tbRuDSxIbySiAwCEcKctpIqpOxoU6RmfkgoNuAixn85A4OSjqFBWyMOl3
39ffb1aNLyQbR5L9TPlwiY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA4IAEuMZf7zdkmNR3LHQU29ssE4/0/N3UAbqpQSPKqXekf8+lU9eVNl+GQ9J7Pi9i
5y+lHQbUbWrdEx3ck1ijKo+1qBcurW0bg0sSG8kogMA8VXvZ6b9S00xxEYIKU6L95NbTQbZbjeninh5R3MQc0j5O57mxJd67vjAmlszD9zd9l4uPSZ4zoH2nlxmUWHNo
L6JtsP01a7+yjs8x2wDQnKeEgzPHDczuKmbNWWK2hrau3hYx+Wza/QhHqVpuS4SXXxvl1LH5DYyIN5cZP2LRh58JQHv+Fl8vPlgIggkA2of0ajALVTE0BLv5Cjf36jD6
6UwUkctWWtQZvGUpGT04DkaWodjovdV9HirnIMliE+ti103NsSyFzvlHYsZocqlbqp4B/AU2ugmS++1XtXSX7V3tJwDxg01Z8aqOVt72SgbUgD6DYOP4ENGX+nf8mvV2
R32tvGDMbA7MsG+El5jMSL5y8b7qqMxZZkrBAlpUqiEl3XKDrrZCZs2+nOhVhkq/mjNViz7s+zAGwKjznFgswlsGCMs+e/luSh9gCz05Jtwp2gI/T+aoid7RNl68x2qf
MXelSorXtr3zdFgo3nwtaPvFslGEU7IMtrk/49KntrvHT2MRBrHpvHAL1g3b8OfAnRu+6k9KS/9uQT10PQ6gcuPFX/ktc6W8DwRNY1EYffn76jB0XKTasgRWOT9xOXA1
iYSVv8e4cn2QMDOmaQPOk0FgTrubRonJFKmVBt0hleoIFrsHzk3H7lCvelokb6NPwm/8zmPnyoypzGsek4eSXJjHNdew2UKnhvAenqR6S8Kcfu3vj+HhdKs/Jsgv7+8t
QaMsOxjy/GPl10nK7l5VRVQfSdeYKEwD7vSA5VpByNJibuDieN6/6YLGJ2h3d8yS4dhl2diLTXpjix/DfNxvPBLJscF3QF5S9Tc1gT6HWFxAVbqGjBe2Zdx0ujOugh4V
KDMz4QixNF6Qxsd/hzAEn39V5lnijLjFn4O8rkIRQ2T24IiVtviTcseE6wqcc8mcX0j36mGKvzWeL9/2+t1qa1iiM/UPb8MeEeONk3N2ya+KntN1EFSRi1lI9KPESs9l
6F4s43udAEC7Ewdf4ATS6AHE7xfIMKKDCpigK7+ZtPCkP6Ul3cGX1td93WzKZOsEiWAtes8YLIyPCQyyEKubnlWECSNLviN88Fll/egmTNTcQAB634fPYac6XOagnjIZ
/wCw8Z9KwwNpYlpQeXe/v0tAniX4fmXQFwhR+QEBzWQhouFBjQEC0ivU3mJhfhSE2/bKtlshAIdjfLyduhFtRs2aMlNcDyFQuiZryB0p1A/K+iJcj8DOElRpZVWgmqGz
h9Z+XAjvF9XWC2hzF6pcYnTOw2bC5uqwslyHThTSYDlbNdTc9rMOwrISgUhPI8XqkiblOP8e/RSmtzq3Wf7EikCfpz7gPlMGrkvMCt9xBMeaIj3frYsws81ln2baUsNG
u2bKwWj/Z1yRaOVbk4VLPa7eFjH5bNr9CEepWm5LhJdfG+XUsfkNjIg3lxk/YtGHdXuy/IyEY72CUA8vkB7YudGWBnod7x8eRXeOfivovXNi103NsSyFzvlHYsZocqlb
pfzyk3jOCV8dxFanDmkhM13tJwDxg01Z8aqOVt72SgbUgD6DYOP4ENGX+nf8mvV2MGMS4Xx329ujW0SCvTu4qrPqzge+g22Bp+dJaQJvBsD/2KgJoCR8U1cLRzF4n4Ur
NCvsqNaJcnmTYbaXAhR8j7qouqUT/OGxCueoits1JbGOz0jFeoLmNVBTovuV0iaNdJALm99oJlbWIUAK7CpzmHO0HApBcsOHQy/RJdkUdvbaVKbbzyLxcAKtOPt6xhTK
YdoHO3hryDLfVbG+6EzPQaqWofWQej42EznBWgiReSCiqoFxbtvB4uLGPs4fledA961Kjjok0iHYUyDIOR1YriGmoQYY4gBbnZzkIC7o/ZTAQHC49OuaxebJZkWhm7dr
BoQjQa6P9UL/OxmALlRHDVgVgjvMnXvXQAoVMBMriO7xvSqpKMYOBxXvuIPGZSx0c0DQvjIuMXiDEwmpKy+tPQrrn5tQhV/3fyFggDdX601c87IOTcgLSaToZt+lYHjU
tEF1ZNnl/2GbaHRLrwdo4bBroL4L2GrfpRyP98djX8kVxXbHaM/eHh5B/25CWXlHAQ5cwkIwxXIfEoTaqduFWalbnXuGFUUmtV1GPME/NEDf+Mh0/le99n4WTyi1qbd+
8zCgmQ0LWexoeUHeJEUjZ4vv+0sdQ9IRSSIe0MBUl3tETAemUiMgBbUUAAK6QXzX2mZRGOiK6qjt2jkWinUYR/wK8Uv2deupdm8CKghvT/toNgucmuqq9EK4s+ft78Zt
IEKzspnAt8XBHzDV3rxLdlsGCMs+e/luSh9gCz05Jtxf7wmPjQtLp68J2FQXVc0qMXelSorXtr3zdFgo3nwtaPvFslGEU7IMtrk/49Kntruyly2BmVn0j5C/9xHXzZAi
nRu+6k9KS/9uQT10PQ6gcmQj0fd6OBNhkJUI4vKovof76jB0XKTasgRWOT9xOXA1iYSVv8e4cn2QMDOmaQPOkwxLdj+IJ7VIY1hz5JDjyukIFrsHzk3H7lCvelokb6NP
wm/8zmPnyoypzGsek4eSXB3EYrkCJU8opuNyttaPnwicfu3vj+HhdKs/Jsgv7+8tQaMsOxjy/GPl10nK7l5VRWmelcic9MgtfGGevFrbgLlibuDieN6/6YLGJ2h3d8yS
m3V/5a7xPZ/gTzeEOhDsahLJscF3QF5S9Tc1gT6HWFxAVbqGjBe2Zdx0ujOugh4VGli0UfmptFgHU2Hh7aiRD39V5lnijLjFn4O8rkIRQ2T24IiVtviTcseE6wqcc8mc
MqwVNPiegNWLxvotwD+eZFiiM/UPb8MeEeONk3N2ya+KntN1EFSRi1lI9KPESs9lypv0KUKQYRzxKRvQ8HzqiQHE7xfIMKKDCpigK7+ZtPBakz5mA9SwWhVE4udfYGEM
iWAtes8YLIyPCQyyEKubnlWECSNLviN88Fll/egmTNSucR/dkfXqWBZIKZ4oWlCD/wCw8Z9KwwNpYlpQeXe/v/Gtp8ctEDHkZu26+yQoELIhouFBjQEC0ivU3mJhfhSE
2/bKtlshAIdjfLyduhFtRk/2EYPXJZ/zn9he4OVyUI3K+iJcj8DOElRpZVWgmqGzXuSHOuptFkGZ3PUZV6lFx/xDDOtOocAsoPaAKMPueX68jop5aW/COGtJqwFsPwVj
YdoHO3hryDLfVbG+6EzPQaqWofWQej42EznBWgiReSCQzFz6gnnm6+P3hM2kGmFD961Kjjok0iHYUyDIOR1Yrj8wNNkjyrIlZyuCHKsqiBfjTIiQpk8hbl3MnAKu3HaR
012N3uHPb6S3R5851LBilaVMDqoraDZ71Kb5Izgx7dtwNQGimAJpBpZ44D3HVtz0BVVQtetc8YoIQ8i21+w0MsbWWECEvNmdebovpWQPdMOK/WfA5bsLNwvkQGte8Q4T
wEBwuPTrmsXmyWZFoZu3a5Im5Tj/Hv0Uprc6t1n+xIpBfVny+0RNFGbfX1OdhB7aYm7g4njev+mCxidod3fMkk8GfWOxq1Ln1DY0iMaeXcwoweOW6R1DOJVvWHNvcmKB
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAQZOdhesV1wK6Vvh37Gv54TMQ/tSUvRznPeVV3XOEC6GPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAP+uF6g+zupS7YGw5830MWHLoaN7lt6s7BsOcjXSBAs1jDimA85Y49OwF1Q61Tw+R
oedhNyJ4AU4LhBzwlNF9D4+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMByWpPySHIVOR3OS7Pq7lrS
Ztq4slqSb3rP0KJuhjzm/4+1qBcurW0bg0sSG8kogMCyg7K+KCsoLW4Os6mfpwbAXMjtqskOS+mMwuHlew78fTmPx6tF/w77VbvXQVm3gh2PtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwM5aJJGd20h6MHIlsPuJ1T9vXFoUdIR2WgoK0xeJll5U96oJbOfj1ameJnRX2AoCpP4oT+UN1Dw9JoPClx3To30iW8dNu1L8uYnO3Dvob4Og
Cn+06LIwMjX2SUnPhoVaQY+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0/srX5ukmawO9lnRLLGOex887ANVgrR6o38OFKio/DKkKSc7qr8MB1M1Zc9QIS5HA
j7WoFy6tbRuDSxIbySiAwONMeHyLPjBXr+vDz9vDfz/nZGmMth7b9yUhzLoTdf3FxwYX05P9R75COiSUkkR2bUal4qu2bz2U8SsAXMNIsYok+LhDiIuribfZmvWmKpsG
fP4TWNHH1O6fuhEshCZONqnpMn9pbePukKjiwmr/HYquyqK5zsQU91e38KhTvTTNj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
FxaqimBX5JGpLvbDnFM53n+POFkt9tftH2bNuXxh3GCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAUKCn2/qSdR0lHSaOSgLLl
T+sMHpglTNq+ECLAJvAnaTozyVMUvslFmyESjTSWFDhVpU3V3m1DSETr6GkxzZTks8J2fmX4jlMjDdAa8mN+Fo+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwJUqVCNYvATBgTHam5A6It+NHKZcU/sIHLJjMNQzOmt7j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAOJeNJZZNPvfoOAGtB8cJW
Nnclnn3l6bYqtSQLxxce5lcQrjKoIilvjhKDdDWGMmmPtagXLq1tG4NLEhvJKIDAzM4nXcdE6ECvYzuMWziVIcbKCGBuOnXLvRf+TX/lDmtxACFwVWGawDfOxMlmbwXj
OkhpvZ3nOhl1iBP1R8GRVnwOqfmbWJhiY3w3ECndOMQOzV0G+Di1WAydD8ihz9O8CecJlBlw60XkxHjp3syWbVx9pa7XSo2w7Gj5lRIp8rnB7C+adtfrbUXq2UK9otwV
ti7reUJd6PADKKs96ybsuLe9NoFAywntTLQKnyG+C9uPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwAEWDk3IDWaXIxoo5gkKK8AqRo344TDG8+HZ7ldtDfnn
jbh8m8wglY279BkklmeEAI+1qBcurW0bg0sSG8kogMA8VXvZ6b9S00xxEYIKU6L9CYCk7T+q/D6jHzyJZ7mopyhT4m5tqx9cgrbqf3I6UV43FPSgNEy2wanKbrdym5FS
exYx2YYG3WGL/CLU41+3vWHaBzt4a8gy31WxvuhMz0GsO31u4pXwIufUYcjdqtbwWfOI1WPK8o6JxZ7XEpFOYAGDdnTA1Jy2cbM2CaFH4AWcfu3vj+HhdKs/Jsgv7+8t
gsAyfx4lTl2irQf8onIoYjxB/4ihbLgIpla94a+bjlQBxO8XyDCigwqYoCu/mbTwkjYj+ZupqEUGyxSMjlIkpWHaBzt4a8gy31WxvuhMz0HeyCOIPkML9N8CiSvpZ4bE
FPz8aXczoOiS6La8qe37ERXFdsdoz94eHkH/bkJZeUdpfVdIm20TU9sC7v7IRWTqutLk5ByMEQ6NrzWK/MBIieqyx9RjHA3VyymhXIhIfSlh2gc7eGvIMt9Vsb7oTM9B
YCxtfF/7HjENRPlP9x1ohiKI132uoqmFU61Au5XCcOsE0wqO8pVtq2XfXadFD4R3Xe0nAPGDTVnxqo5W3vZKBrRBR+kslc6pQPpDoRhc6764dDZ1Q54pa0HcFjnLK8T1
961Kjjok0iHYUyDIOR1YrkvHzBbmplGJxe4xhh4uqJGcfu3vj+HhdKs/Jsgv7+8ttHhSZNnF95lrilz3SgaL1VK6MioFtVE5tDPCjz25oTgBxO8XyDCigwqYoCu/mbTw
iv1nwOW7CzcL5EBrXvEOE8BAcLj065rF5slmRaGbt2tMHHo6I3/m0eiVQe4c5DZGrGrZMZHXxZavxEInMwfgZd7II4g+Qwv03wKJK+lnhsQU/PxpdzOg6JLotryp7fsR
N6Ze53psYakr4J6/5Dmlh1A10rv8WA5cmVUG9ZiEp1yPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAUKCn2/qSdR0lHSaOSgLLl
PpiLbDw4sAfC7pWsCXv4ANUl80iyti98ZcxAanPdbP6PtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAvvWIIJanZhqLlJt2oDeHC
hnKU53E3ivtTsC+q0aEVsZP5SHbn0XXz2m5ZyW0q56GmS9S3uuWbT8Yk+wl/cXKY2HPwHnLWyOqANJfdiTcdhY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwL3v7twNGVDoDtpQBVOA3r0+lMR0nSm/Kgsl2p+sB3/qj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMABFg5NyA1mlyMaKOYJCivA
TYDYVpgKKzkEXXJpb5lXzI24fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDAPFV72em/UtNMcRGCClOi/d4LIMiyjRsm8pEY3KGaXm98q7V6DhvySELVYoYu0KZZ
1Cgwn84sWISzzS7FodDuDHrAtGIvbA1Tj8UcDVNoL4RbNdTc9rMOwrISgUhPI8Xqc4P2kONHgqskGsQRo59xxY+1qBcurW0bg0sSG8kogMC74w4wEBAepOCiQ0nq3dzK
yNqhAmGR66FlC/7IqUGi3d/X329WjS8kG0eS/Uz5cImPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwOJ5/HIckCv+0qVjtBIomoWtHGEH389Yt46KgEw0U+WN
uIEbXqUhMmSOjb5x8EaeF8OFqSHF0Hmjrcs0rJIdlFNkaewk3l1NwKwJ0+iTvk7iC5rNv5YNh+dQrolpVWpxj5X7PY7C1VOuy5A6OFKGQsOPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAsUofP4oR+mub8YV8qkNomiTCEhsuPlZc7SUC/zoy9mN+9BgSs3/5rMjuVLkIHYQT
O37HJSohuWa6bwgXSytYmpry7CZno6e7msbSbDsHpiwBDDpy8ZxVwIZ4R1oZ2qPSvRpidAjjyVBNWuossTi1d0lzNguq292MFFjOH1fCykJctbZhr8mO8rvDpluOAknY
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCcb3dPwvsvcvwJQW9sFxss6AwMMCcY8oLmkEVIF0RtySdCtfuGIUam17WdlqxVEZCPtagXLq1tG4NLEhvJKIDA
L71iCCWp2Yai5SbdqA3hwmwmOnctcedKo9r0lP6ZqTht9WViA8WmJZvLmohu04WXMXelSorXtr3zdFgo3nwtaCxmJjCXxdxbAUg9Aaijw1vwfrCRptDZY7a77CrMRke9
QOmdxd1xdmuYTZ+769sz5ilBdl+9IAd24G+umImQqqtWguVr0nEhmMg/uPwYl4URqSZ3kT9vKMpirinOSr3oFL04RagGRuK+RHdK13JTEEez6s4HvoNtgafnSWkCbwbA
UL7dXYAZGv9dwYRlTqGSAgpJzuqvwwHUzVlz1AhLkcCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMD4d8UZOOKLnVTEyU/ivuJG
y6noOc2/5n7DanUKahvz3bQjDw9WQjnAG9HtFN9i94+PtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAvvWIIJanZhqLlJt2oDeHC
hnKU53E3ivtTsC+q0aEVsZP5SHbn0XXz2m5ZyW0q56HbMC3eKPRRWGKNFJtivHq1VU6gyGuofmgxly0kXAaY9I+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwBQoKfb+pJ1HSUdJo5KAsuXal0mJcmVfwtQayTibYugqCknO6q/DAdTNWXPUCEuRwI+1qBcurW0bg0sSG8kogMCUyKszPv7Goe8Dl/1zunss
6AwMMCcY8oLmkEVIF0RtySdCtfuGIUam17WdlqxVEZCPtagXLq1tG4NLEhvJKIDAL71iCCWp2Yai5SbdqA3hws4IgTMlzaLDyGTCTaGNGmhuD/GmeI5gdpp8K2wuO9Cx
SI0hdsRexE3+4k9scLAzqPa4hB+58ToJw4P5oqI7WLmv/LNXTuPSYDIw9G+vPslfLZJCROpEA8RwIbZ+YOw0tY+1qBcurW0bg0sSG8kogMAUKCn2/qSdR0lHSaOSgLLl
3sBlj5Qea6d/wgp0s0XRr5h2dpQj3fWEEJKcOsOi118oweOW6R1DOJVvWHNvcmKBj7WoFy6tbRuDSxIbySiAwPMFzS0KwpEVQkOn0lQ/es+Ka2sPZpMAoe0GLGjgS8V+
S87FriQis0GeiGcI6RGduZKLSWABE75EjF4TcmE3p0V3MNfjRAgvUfHPCvcidWKfiWAtes8YLIyPCQyyEKubnqczEBQRlXtBakDPuOtSaWd5XqzUaPenYV857XqC9z2h
oC+E5Dsy0uOcDbYup13CnqLOUei1EL85J7jGNvcxf7WPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwKEFiBwQ4AvPApELb9S857rl9O5ISnnwi1qzxjj6IM97
i2jjPF9b9F/yY+yGZnP9r4+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKDMXelSorXtr3zdFgo3nwtaNaA0B1mfrWTOSMTmfmTv26Ac+ph2ckLpS3CD/1GIUyD
izJtzE9mSYn500wjm4cIIOGhOJYTLKOdO2SBMHMp3HBd7ScA8YNNWfGqjlbe9koGpGbGGi2sGgZgpcoLmLAtzovH9BXI9w47FB3KaqIVq/tibuDieN6/6YLGJ2h3d8yS
iaTzlaPCnc40cMwdpVVH++gFx940ioMN6EVYCu7qiHyWqZem/kdbUiAt8L7aFRP4EsmxwXdAXlL1NzWBPodYXDoLgiWygBgWyBHfx7/Y039nWhAyGp56Mn+Y+XL/+KQR
8b0qqSjGDgcV77iDxmUsdJoiPd+tizCzzWWfZtpSw0bRT18AuXhpkRPjd77EtOJBc4P2kONHgqskGsQRo59xxY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwM+jeqLf7F0hlf3sATGgk4QovSmQZMfdSqD+uygHVRBujbh8m8wglY279BkklmeEAI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwAaDiVsCDvQgwfmHf0imfy7dxvKh9ZMhw/36feIv7oOk8k/h8VLp6SKiwk3B4VW6gvK7ye31LpLAcvvAp5j27Vdzg/aQ40eCqyQaxBGjn3HF
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAYzo7S+/XGUYuj9JQn3nuYy9TC+PVR7Ebe+C8+bq23EGPtagXLq1tG4NLEhvJKIDA
Hj7F3Rz6xogmkhI/T6QCNP7K1+bpJmsDvZZ0Syxjnsd63xvi6GlEUJknxEfSAgvtCknO6q/DAdTNWXPUCEuRwI+1qBcurW0bg0sSG8kogMBKYTRDgMVBJHeNlvVYNYl9
Y9uALeCxzMSn8ImNa8s3tYkqX88ZB7Bjb1HxD29Obrj2Vcj+jiwOEk1QU3ve+XbIuY6qnH1KpGVFJ30BNN/dFLtJZnqwgRhB0ICyvybncy2uyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwFSGVDqrFDOKMvWAxSKFwf//2fndZGf7QBiHh3FLsyphLZJCROpEA8RwIbZ+YOw0tY+1qBcurW0bg0sSG8kogMAUKCn2/qSdR0lHSaOSgLLl
Xe0nAPGDTVnxqo5W3vZKBq149U64o97nwEyakEtakdzOLV7GN3no0Al58AhQvqGQ73dPnyWAlBZ6BLQPC1ej7O3+qOHn8Jd/LDNR0g1h5SpYojP1D2/DHhHjjZNzdsmv
kmftnkEWlhylnWhWpRijXeckAVFMBTXuR8s9QTXd9HJUnsRlrmp888RxDgLj7QZrnH7t74/h4XSrPybIL+/vLXOD9pDjR4KrJBrEEaOfccWPtagXLq1tG4NLEhvJKIDA
/+wzxsQVeOYclHF8A8sJjBEItNnHk1ciFYqm9DDw6/1m11TjRVgCBvAXOxUjeWYRj7WoFy6tbRuDSxIbySiAwB4+xd0c+saIJpISP0+kAjSwY/brEb3Yv/rAKBS1bNvh
l+m5+reZ17elfNL5MAkvCtf3uCY4PnxZRg+EKc5pn3Kg1FjjWnqYbsNXT6+lEW4uWUvyt6c3Z1V9R2Aqb/hR7vC1mfe9QBWZxeYbkMsftY3F2h0B2deyhZ9l15iUaTvW
8RIDMX1WIzTaaO4sNNC7PFD6+9P37fshasBXyzTW1Cto2MXqxCsCZNX8MXsDFsHASsTqh79Y6LTORyw2PhIY2AluwhJvlvl+UEsCvFijnfZxoc5GcP2CLHy8qP6Ib5Qz
Fk09tdxPxKz7DkfOF1A8qtA0pAVbV4BULcYXKoWJBFAQXo3+wTyO+HudCMiaPfi0lQzcGwv6/QNCDqhhgIXe30xAUUdAwmH5KNoMfp98lh0JIIfeuDH3d6EvRvdRnNsu
OTvqvI7Ihg8NR/E+GFxcokadhEPByXnMJ/5tj/wP0oLRuze7KE8ld9XhJWCImbjI64ViDcPbPvf21TJIQnYjYB+CrboySRGCKsvLy7JTa0TKBtg6Vv9lgrc3nm7u79ii
/PCe06OLkw3hNsf3VKBKMr55sBDHZfokV+YUe9o6uEgZTgaROR465PklzJcOgKBsMXelSorXtr3zdFgo3nwtaGNTzuU1npxzz6+k3EzQeW0jMeXwrwUm9EeGeZU9oPTr
961Kjjok0iHYUyDIOR1YribyyQ+TYC8XRWS/0KrpcgFa1kUq6y/EN54BtVRFUPoKjun0GM9oFlf1b4FJVx4C3mSRyQ28jUKMHtn3x7Skuiu5zrBJK5PDCjPWkpEUTwHh
bbveRSnRu1owMGmsszz+2ZblMXpMVNAFLmYomUeqWS7pm1fRX8xRAjSnaC8BgqiFAXV0vr7Vflid/jydETTQ6D+DKz/4CUAhO8tILumpFZTFW1ag2MWZ4qcu84DNWsi3
XtwSmXBlwUpfL8sTS25nYOPWydXcLhQWPLjm6ppBxqdJld1HA3ixoQP+zzXD+t1MjjBQ75PEGCAZy4xAQPPuZ3d1IRVmXDGWZMfVRPpnWEaglWpqJYb3/7jPXa8MxJDl
Sv8I3Yzfygc7bJ/prebLZ5QXQb7ExWMx4KPruolrI1XioFpBX3YvmfTdMzYpQveg+2uw1C+nx5o8xMhYcjWmiobIyJBBNlllJLKpMqQUQ7TvwGoxOohuVsfcz019J0S4
SZXdRwN4saED/s81w/rdTL39waq32F+WvvrV5SeID4NDlKvfSZvKB8TAhOUgh9xJJt76ZC2HhU3koN1eDD6Y0+bxer55WoY0JpEvL4ySUZOXwRD0+9IVJ1Jaiyr/s+x3
353KcWcYd0YIxHhleFffE20GuhTb7qMiEWYCUvCELo5o2MXqxCsCZNX8MXsDFsHAjY7GPPaHK8+tphsjiY08Vy1XdbVlel6dVRDXRZug6kRc87IOTcgLSaToZt+lYHjU
e9jlbjMrvwel1nnwARX3m9GWBnod7x8eRXeOfivovXM3vjQTRayQ8EyhYpxyBbRYz3X0LoV3Rp/f+yAQ34n7iq/3uA6It9XuAR9HE2bPexOPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAkN4g7GtulQm4u6gVYsLh3wv06vwl5vrjn38efVSoRRCsHdT1W64HgIfzpxQSxSymx4nlgV2LHX99jiDVwF1oD
XtaYScI0FKTU6fAO4ILUEOZmBZuDE0NVHfR3zN/xZMKPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAvvWIIJanZhqLlJt2oDeHC
hnKU53E3ivtTsC+q0aEVsZP5SHbn0XXz2m5ZyW0q56HdjyT592Msmc70Bpa2glHxs8J2fmX4jlMjDdAa8mN+Fo+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwJUqVCNYvATBgTHam5A6It+NHKZcU/sIHLJjMNQzOmt7j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAOJeNJZZNPvfoOAGtB8cJW
Nnclnn3l6bYqtSQLxxce5lcQrjKoIilvjhKDdDWGMmmPtagXLq1tG4NLEhvJKIDAzM4nXcdE6ECvYzuMWziVIa0aXLHKMNgqmC9emQE+o3U7VTE0pXnEDNPPnEnTgYDN
hGl9k1gnP+AtJSn3SwPwphRFxbHU2DDF3J1Vsblaic1m2riyWpJves/Qom6GPOb/j7WoFy6tbRuDSxIbySiAwLKDsr4oKygtbg6zqZ+nBsCl4FrruIwp1LZdANrwJGwP
cIl8IpNngRSwfGM/X2Q0CI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAzlokkZ3bSHowciWw+4nVP1pS8Tk0b1tXZFEsF0Ds5YGo/0aalXpaG3yT1tlKazuf
wtEh1Cu+1rU1oWFiFoj0Lbl2OpNH7RlLe9O/3HN8IkL3g1EjwuxZ/dRw+AJv1Krf+cRFthcqO0zhhSoouLurNCLrFZE5mDrON2bepVGaZS46FE9NYqGj1byqo/zRsKd8
U6ykRv64vZNyYVWH2xYxA7LgrjxV+9kQfdyfsR43wRQJg/p2vH3DyP67lAndKoZgNQpVqKr1ut9h34wvesr5Ig/k8cnEVIEJld476lyT25QfG713j092A1lDDCoCTYXX
iWAtes8YLIyPCQyyEKubnibNnWGlRU+/IPTeQ22Vozdn+uGBBbwKI9GSXdxHT3TKNY0GNernjXZvN6v3mzUaFbDD0OF9Wjru9mQlfyTfdXu5GIBgOdHnOIlmY8M4RICE
sEqGr5FwNzh2VRv7OHmwm9doEkHUjx4VSegb009vl1FvhM4mCt9Swc8rsQ2zBIIvYm7g4njev+mCxidod3fMkk8GfWOxq1Ln1DY0iMaeXcwoweOW6R1DOJVvWHNvcmKB
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAt+QyWL9P+3AKQi6ACI8HAI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMA/64XqD7O6lLtgbDnzfQxYcuho3uW3qzsGw5yNdIECzT+UD/3kJ/dFH0UmPnB4Q8QORgc/PE13P3Nu+K4ZNaUS
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwHJak/JIchU5Hc5Ls+ruWtJm2riyWpJves/Qom6GPOb/
j7WoFy6tbRuDSxIbySiAwLKDsr4oKygtbg6zqZ+nBsBcyO2qyQ5L6YzC4eV7Dvx9OY/Hq0X/DvtVu9dBWbeCHY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
zlokkZ3bSHowciWw+4nVP3il7fBGzy9JgcZAlvUAkNACaddhJMzOW2VWv5kutnud9aTmMc5RWGxiQupxHRo8Go24fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDA
Wf5s0PuxtgTUL8+pRYJYzl+7inNcBHd6gN6BPholOU2vC8UpWsZhE6c333ksRUwuj7WoFy6tbRuDSxIbySiAwIkTtD4+JQAJdIisJ02TW4xbNdTc9rMOwrISgUhPI8Xq
6q+jpzuIsEGRsfUsB4fyY0y4f0mgMwOlhJWN08Ud6bycfu3vj+HhdKs/Jsgv7+8t2Sc7Zhd9KcodkxXxihridYhWMtCc5CI7xLPt2JCfx5x4zPp0v7BakU4coK2FswLb
MXelSorXtr3zdFgo3nwtaP4z/6CdUx8SrBA3W6OjUCrSYa84rBfOxf8202DjTenas+rOB76DbYGn50lpAm8GwPOKgXnvsOOIO0lzwWAbqIth2gc7eGvIMt9Vsb7oTM9B
HqvN1xLeY7McMISjlUqBPHl6yzhVLlcXtxiohkB0h/MBxO8XyDCigwqYoCu/mbTwWjLFV852TmX4leCo94HFXKlbnXuGFUUmtV1GPME/NED+M/+gnVMfEqwQN1ujo1Aq
B8jhBPzRrGjpQlaotBzfB6AvhOQ7MtLjnA22Lqddwp5fs4LV/cQ2Zgl8NzxSMtFjj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwFLTH+Cju89gmooP9uGI0je7isQz35ZSCeivG+BQtbsMzGf8LGAR0w5iy8v80W6UuI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwB4+xd0c+saIJpISP0+kAjQ44cnmxCQanhzaT2rpViJaDd02YRwbKk6Sr0qhwPhOk2My4K+JuKJrB3kIDBj1sP+Q6pN/9vVEfjV+Gb7SVm35
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAiRO0Pj4lAAl0iKwnTZNbjDz6HD4704TGLdc87nXo1xFzg/aQ40eCqyQaxBGjn3HF
j7WoFy6tbRuDSxIbySiAwLvjDjAQEB6k4KJDSerd3MqQMetHRbdrVS/0au/fjdxEgNrgm2DbeiZzMdQsWOxeC4+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0
MXelSorXtr3zdFgo3nwtaOaNPBFAwpydRU0W0X2LKn/jmY5bsRcpy/WvGPLSywy+GCK0X8jyp2oAgGeitae54QpJzuqvwwHUzVlz1AhLkcCPtagXLq1tG4NLEhvJKIDA
lMirMz7+xqHvA5f9c7p7LFGmsJbPzdtSR6WR8las0GwnQrX7hiFGpte1nZasVRGQj7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cJdPC2/E6r6xENby/8VoBQD
P2HvyzeKpn4nsA5ieUADJyfEI99GFiw4l613rQBdV0iBbxOgcJp9T8qSfJayiP2bWzXU3PazDsKyEoFITyPF6mQ80AYGhPb2ZAhzDCYxYQ5OvLuwmSE8Kimg0NS/4kll
oC+E5Dsy0uOcDbYup13CnuPhpxXsgMwTBI1O9ITxNoMaSBBgORJvYfnbvAyGWww5uvqkYxGMMpz24cZ+WtuzSgrv4EmzL6OEWroRBZk1Div3/QpkknvDccn+4ix/gNmw
gHCgrqavwfuJtV9/06iTcL55sBDHZfokV+YUe9o6uEh9P5MxkWvfgHasOUhwo1nhCUcdQWpZXcaNeSC8R6xBsUsgybM3850BxNR/nlI77O2QGcAIDoyRJ7aAs0uXorWm
nRu+6k9KS/9uQT10PQ6gcpdEeeQD3ZVYPa7qcgT255+x9yJ/OkdTJ8zt9j+ry80CjzG/jFzq+Pn1HZbuVE7XnX1nKN6LvB/9R6FtJisJJI6aLeVKkOCkCwDHBeWPhsYC
KUtt0vosEMs1TBfpsmupCQDbKx5pdqhVTAEgyIkfIkIhdCQtiAVVWrhp1evTOFUY0BI+jFWwzzciQmAytiF93hARhPQfrhnhnySqcXIXv4BbYaN/ysos1/WDVCBOMLlW
RVQ6cmQus6NHdz1c2P4AFgn6RPVOslEMA3Oa8pQa9eHb9sq2WyEAh2N8vJ26EW1G5o08EUDCnJ1FTRbRfYsqf/A73qs8BC3OcD/K/H6t3v0BxO8XyDCigwqYoCu/mbTw
kjYj+ZupqEUGyxSMjlIkpWHaBzt4a8gy31WxvuhMz0ELLzjvAKlW2JNhw6bBN0UloqJlzws/47enKua+1oVENJoMMLOswX9nR+I8sSsO/wxgSW7TWCcd5YRPQitqScc8
fel/4106ZSkzsy/B+xi8Xr1BNCEogT9mrmgt8mOeZTKiWjCG85FOAxo4Mhr5jDxM8nBuNqCISf2PHR7lDikcS7IZBgSp7oRMJni1Fkdo3i9pAX9RL4e9jMxtIxnKspvZ
wEBwuPTrmsXmyWZFoZu3a0bmmiT18cnFtiXxCvkyKu+Cl6MF9G3hEEY+3Uft1hVUGfC67g2re/wz2ES2d6FppAHE7xfIMKKDCpigK7+ZtPBewXYovg+bEQHaSR5Gr4LT
y3cgMLcOtnd2t/MFKQoQb/HYx+Y9GMW9CcBpcGSiFNVctMg1TXzsB81RWnMyl5ZDAraCG6rOiVuo0XAAE3BMHrJBaTvDcjLXr9uHnU+Tc1DiGoRoW7Y/aBv3Mdtwcyqj
nRu+6k9KS/9uQT10PQ6gcp0bvupPSkv/bkE9dD0OoHKgL4TkOzLS45wNti6nXcKeJqEjyaQSnbH47JQ9W/F+8WHyX3w9WDTEk+GlvhSk/cLTd4qv+pc6MEHpz0YQn2tg
DHTbFXMoOoJjpoaV/N8oo09jg7L/ozaNJkYuB6Sc0h5c87IOTcgLSaToZt+lYHjUpNyTU2FSdsJOS88jgsmByjy08sWzRM9aXnRZCt30/4aRsMINou/MWOYA0M1lEb12
CuFrM2oCKC11GaXCBUynym273kUp0btaMDBprLM8/tlucrm08HmCXWnc8G23L6Kiv7equXd7E2uiGGECCVMGhilLbdL6LBDLNUwX6bJrqQnV0F/8aERjW5pyaKuDBR31
1d6JlEeD2G6sNbXIQ5zFFalbnXuGFUUmtV1GPME/NECwY3mH89WM7ZsiJEuzBovmzi+2QyQ0EQAF0Z7yQInHUrwV3TZ8UPv2c4JAW6MebFGg96O5ZNtO+Zr0ePRhXDnp
TdCGp/P5V++U52mzCbKBTO8otwDb1bplzOQsEclONDV+f7iB/EE1ciyy3ClJ9F05NCvsqNaJcnmTYbaXAhR8j44wUO+TxBggGcuMQEDz7mfzcpr+Bm4Opex8JpI7yHcI
9YYnaeluhlv3mox4AOuS62Ju4OJ43r/pgsYnaHd3zJJibuDieN6/6YLGJ2h3d8yS84qBee+w44g7SXPBYBuoi13tJwDxg01Z8aqOVt72Sgb9vxTA0nhv8yoo5NkofAJC
pGcM0tZ5YKO/el615sZf4T89VFiVld1/OtDH0tIjJaNjch5fTEgBy3cL478npottvCm+b3sEfaZ0lQE5jR3/XnS+/hyH8aLnjf2A161DSDuPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAvvWIIJanZhqLlJt2oDeHCipH2XERREhMosdpriWb7UCpKyE2Y/UHMW8O24j7VLUuPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA5SiUrRk2GRx4b5de4MEhFb6daZ3NqFdCIXDvFOX8f4OMsJ9FjruegfjkJjtV7NQB
qrsfuq70EC0XJBHg9AeiHJANAOUCf7afPJ7OoOD7o6syI1jO2Ge1vybWE8jVlJxR9lUG7U7vQI+SgbT5mPfC5OjxqnxUCBPufEkWou0wXfBwQanz/eeGJUdc0tgOu3gI
qARxq+OVi+P1Jvlvik0x3Xg4aYt8mzERDgnNz2h8e9eVkA8xS7aEOc9xRpCg/IsFrd7zyRsH/IIldsAWYA1k8SazbDdahp4b9PKYF74qCJTX3ZLE1HF61QAi6lAkLWt9
CQLEu9H+awSI8bOeVH3O1FgeUtzxnC1dwYORudv4GQIN6eip9RyDwM/36FLiY3AClmkeE1rZep+fYrWxF1Fst2FX11jpJ7Ixj0iCkdVM+otxgoJ3oRtCtw8bhqgEsHrS
1Nzqy+at10A/iAPMp8YKC3aodIKplYmPQ8yOhWA11rSgCD7cP54wSbiHXrnd1/6QIpoTHBgAOcDmA2ZHR43cqTJvrryEZYDb8NmEvpUCqIZBe6Sf6lmDzmKJlQ6NCs+2
32ouXntBtLDWbvtuoVkX4mTpjY6XmvkN7eILUsJ9w9DnhzvOVqEtFWf4XyIUv0OG94NRI8LsWf3UcPgCb9Sq3/nERbYXKjtM4YUqKLi7qzSQe8atMYx4gFh2KD4yRPwE
9NLIyD0ts1r1PiGbmdkK/ttxEJ3s2ttaqr3Q2Y9DOIDBVQM0Nq2Nuf9vMdjSR8hQUalnQv7US9J5ZdZH07/ZAsWMxll6y+1rQ9ZFa3ytfhYy5iF0thwXMbKbt2cHOyML
0ZeWAvh4fR42aoHWYQQoDsrY7eX/yT/l/TPWlRqLqeePtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMBSJMaqFOQDSY8SpJRSJacp
2+e0IRfJ/+6q7tr9eRuWNo87GyhJeP7JaTTK/C6MnlOPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAZ5oJIosm2oHONobbv/RkE
T7DlCOg6sEXPCMprS2qDwpSRadpOYVFAlOnav3D0TEbRtsBzehe28KeyV5+ebZsOj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwMWoSy11l/ktSZ1vGWfBRaBXEK4yqCIpb44Sg3Q1hjJpj7WoFy6tbRuDSxIbySiAwMzOJ13HROhAr2M7jFs4lSFl/MiX2v4cuhzgzagWuCTu
JMjHbg5sgc5toUk9uRtdVI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAKWhMGB7tD4gfdH++B1seq+yfH1N/tGR7ZcZLOiUpK0p+5no0syJcqgYLCepw2DRz
4Y0dmPFmJatxUQ0Pmomkt6/8s1dO49JgMjD0b68+yV8tkkJE6kQDxHAhtn5g7DS1j7WoFy6tbRuDSxIbySiAwBQoKfb+pJ1HSUdJo5KAsuXewGWPlB5rp3/CCnSzRdGv
mHZ2lCPd9YQQkpw6w6LXXyjB45bpHUM4lW9Yc29yYoGPtagXLq1tG4NLEhvJKIDA8wXNLQrCkRVCQ6fSVD96z6UGtDiaJWtgFHWDwK9MGQBKmy2mo9k1gylffp3+cfZm
EI1+r1EyhwkHbP4Xv1ep2LgJe2WOg69PJ9fu8G4IItOLsBVamRyMVX06Bkd+a4WVj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwOJAHNHtMJratdJ4W9UhLkWWnbRKKkorsNcVdhAXusUWj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwD3fEUD51U89DHJ6WBOKsvT5a2OHWans6c8I0XvaBwNs72D9XSGWkqQYRxzI6zkVsMk/M1183rZai9wXZs3oy/OPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAqMBLf2Y4/l6YixZW9iYGntSMhh79D0qdyQn8MPtk8KuPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAUKCn2/qSdR0lHSaOSgLLlT+sMHpglTNq+ECLAJvAnaTozyVMUvslFmyESjTSWFDi2q6U5cgybzfslKE8jI+J8
s8J2fmX4jlMjDdAa8mN+Fo+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwJUqVCNYvATBgTHam5A6It+NHKZcU/sIHLJjMNQzOmt7
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAOJeNJZZNPvfoOAGtB8cJWNnclnn3l6bYqtSQLxxce5lcQrjKoIilvjhKDdDWGMmmPtagXLq1tG4NLEhvJKIDA
zM4nXcdE6ECvYzuMWziVIVOfMAJi9vhNWRtvnb9QNa1Xgs3MpUltlBCyMDAYTSIUDE/PauHCP2uXs378Oozv3Uw7paTOttWR/ZshRuSM3xDYPnSrlePsUeiJs1pL5b2I
nW6EzGvcaDwOTXKUagO6a1gZrJSHz55DR4lUpvN5TQe3vTaBQMsJ7Uy0Cp8hvgvbj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMABFg5NyA1mlyMaKOYJCivA
KkaN+OEwxvPh2e5XbQ355424fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDAPFV72em/UtNMcRGCClOi/WXSPZ9bKc0KxaEia7CAjTuvg+2/pX6hWjntR/8uDmVv
1apFgyb8GRm15MbgqY4CcCfueNoTBnKkJPZMYQsP+t7AQHC49OuaxebJZkWhm7drWOtyqHuLYqFE5UF7V9TU08Z85gLXbopvGjQ3FkQljxDCuCxbu1g/3dBcZ3tbwN1q
4zmK9H5JqOBS/CDFtABx4DF3pUqK17a983RYKN58LWiaVKvAuqYZq20ypT+/EQj8M96FHz3b0twNbDOzUI6Q/fvqMHRcpNqyBFY5P3E5cDUMSgVP2XUc1b+Fzl5gjJdO
Nxqw1Mrz9DBFgkTXo6pR2MtgNbsRWoCOwMzu7KxXJgQMxIc70JGs1ffk77BfrurfN0o7FCeG4ixkiIMliKY4kMz+LinWhkhYvIoGiuY+sISR0zt5AmR97I6OqtUAzKdD
wEBwuPTrmsXmyWZFoZu3a0CaVCcZfkSHzTpIulaIGd+x7Q7mIFA2vp9hwuQC9LRTTrA8eA4hWAq1K00bUBU8cfG9Kqkoxg4HFe+4g8ZlLHSYY/bUEpAjA4jbK13QXXxx
XLTINU187AfNUVpzMpeWQwK2ghuqzolbqNFwABNwTB7laHtFtJcLgDVGC77uRZXmyqqw23oZiBJ2IMq/JVJOov6Qm4HfEQIwAc/xwkfE/TFibuDieN6/6YLGJ2h3d8yS
ifBsOYHC7REuJipnwHIbY6AT1cAzgZKCfsq2DOr+V9udG77qT0pL/25BPXQ9DqByx4FFOzA0qsZI7IsMmYCSEcqIJtEmvYeBjKtfeWMCbYiAz0xQGT0Cvdq9LLStWkEj
wAKsREO6Zo96UlcD2abCatv2yrZbIQCHY3y8nboRbUZbbYojc8j2vqxEb+qvLYbdhKhhbit87Zr7k8Tdd7kJs2HaBzt4a8gy31WxvuhMz0EXRgYprQ9BKGbOa7s1tXO7
6w81++quB4tzWbKGeL29q3nQkOmrh5Tzr9bTOEU1UMLKiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiPwj32wdQnUZxdDenFIVl240K+yo1olyeZNhtpcCFHyP
jjBQ75PEGCAZy4xAQPPuZ4grPv1vK0/pMVFoZOwRrVVAq9yL6lXFr3i8s6s7UqkJBrCQBzveeJIPfkvgX3gFxlVNwkOh/ot3H9v+frwYjEISybHBd0BeUvU3NYE+h1hc
yogm0Sa9h4GMq195YwJtiNieUvpaF4Z8x45uy6TMjZZnUTyIJH36AMkxBKclh3ozG6FlFZlTLSvAPZpN6SkyTUCaVCcZfkSHzTpIulaIGd9Fz3OyupbXB08jYaKA5ZI+
auQwNP2RRb2b2XJ7gPNUn5oiPd+tizCzzWWfZtpSw0bxMwnCSwDOdR7CjlJLSyEjLonoBVX8ZUJ+nZhayqGyLMBAcLj065rF5slmRaGbt2vKiCbRJr2HgYyrX3ljAm2I
JqfggKkdEPwnDMy5Zoszo5tdJM4WzE+aFtJ9EK4T0OzKiCbRJr2HgYyrX3ljAm2Ix8ouJdQTLlvc/URxRER0w7h0NnVDnilrQdwWOcsrxPX2Dl43NsNYFOrWQkGsrVdK
kz+nwTxmLIydUb4eBQkzhwHE7xfIMKKDCpigK7+ZtPBqK9lkc8hISUDTav6paYNeyogm0Sa9h4GMq195YwJtiMqIJtEmvYeBjKtfeWMCbYiTHXfcvsY/JEJ8v8NU9PCX
nmFo83c8IazQxWNbcd6dvNv2yrZbIQCHY3y8nboRbUaj6gK3qXKwNJSbEnEu9GKpewALxVkfM7TpWFMr3FtnnMqIJtEmvYeBjKtfeWMCbYjNlMPavjZaG8kxX2u8SBTP
rRe3vUroauj4faft9glLsvwK8Uv2deupdm8CKghvT/udxfTHXTVQawvcNfIX4kLl0UKcUnCcuGl2a94ticEHplGgF+1NIXGGc0lV4WreJwbKiCbRJr2HgYyrX3ljAm2I
rLtZ2/GNaoCKtvS4QSQCxlK6MioFtVE5tDPCjz25oThHn22tW9H19vIqo0h599bqjjBQ75PEGCAZy4xAQPPuZ/OKgXnvsOOIO0lzwWAbqItctMg1TXzsB81RWnMyl5ZD
AraCG6rOiVuo0XAAE3BMHmROVRZfkVwhvQbMl4tlzIdiIULQKgKyRypHAaA4theEyogm0Sa9h4GMq195YwJtiInwbDmBwu0RLiYqZ8ByG2NHCnZQmMX4A142F2M5bSoP
yogm0Sa9h4GMq195YwJtiKD3o7lk2075mvR49GFcOemdG77qT0pL/25BPXQ9DqBySSgraxeGkLmwUFDDBc0XlYeeu67xMEuyL4OqH4TMEWDKiCbRJr2HgYyrX3ljAm2I
V+uNhopg1SrJWWrbIBaRno4wUO+TxBggGcuMQEDz7mecfu3vj+HhdKs/Jsgv7+8ta0lOJOLGXKjvHC0ToMIwYRZH49KSWdP0VriMydzUmAnEfaJ0b3YWK7DUKrqlagsP
dLnqKtVTR6FG0FWc8IzPL8qIJtEmvYeBjKtfeWMCbYhh2gc7eGvIMt9Vsb7oTM9BDRwpWjzOkcDgjl1Ws0gv4IT4DVNReH8ZE+rNr6kOFJJPZkHrSd/YpD7yJ+GkWart
yogm0Sa9h4GMq195YwJtiCyGVvHiCDNLQUa2OifRrh4kwq4bH/gFrk4Ru5F3ViWKyogm0Sa9h4GMq195YwJtiBThOEQKZ9IXJ7ZAGgEcrbGQsuoNBMFG2d3S+MfcyTVO
yogm0Sa9h4GMq195YwJtiFiiM/UPb8MeEeONk3N2ya9AmlQnGX5Eh806SLpWiBnfnifbija+sB8ruJRhqSlUlmrkMDT9kUW9m9lye4DzVJ+dxfTHXTVQawvcNfIX4kLl
m5Kz+bwor+x2sxtBTII1to4wUO+TxBggGcuMQEDz7mdibuDieN6/6YLGJ2h3d8yS8b0qqSjGDgcV77iDxmUsdEesNb9RG4BYVf2SWCx4oqZ5UT+z2F6vClbOdAHN+bYe
yogm0Sa9h4GMq195YwJtiAS9adVehTrvwgUg9CnXZUm+H0cKxGie6OhmRPtkysE5qVude4YVRSa1XUY8wT80QIubBCQ7I0hsrM8AlzGtZC5mxlpkD3hPeQFJ5QQ/cndF
XERkKwW5G95ByvbBAuVEYKsukoXo4rMrRUM6WWUw/WqOMFDvk8QYIBnLjEBA8+5nWzXU3PazDsKyEoFITyPF6sqIJtEmvYeBjKtfeWMCbYh9GatTzk6exGHL2TZteO0i
omBEvlr4X1gMbkn53ehXN7wV3TZ8UPv2c4JAW6MebFFkTlUWX5FcIb0GzJeLZcyHpS0qs7mBOJs9DhwDWX64acqIJtEmvYeBjKtfeWMCbYj3rUqOOiTSIdhTIMg5HViu
mGP21BKQIwOI2ytd0F18ccqIJtEmvYeBjKtfeWMCbYgxd6VKite2vfN0WCjefC1oyogm0Sa9h4GMq195YwJtiOVoe0W0lwuANUYLvu5FlebwO96rPAQtznA/yvx+rd79
DRwpWjzOkcDgjl1Ws0gv4KRsgPF5b08WfNlg2/EOGzc5xOEFLHR3e3sufri8tCVJi+/7Sx1D0hFJIh7QwFSXe8qIJtEmvYeBjKtfeWMCbYhiq0ya44oBmX/GToOs6Y0Z
KsSu+sxxy4FvypJS2XJavMqIJtEmvYeBjKtfeWMCbYjKiCbRJr2HgYyrX3ljAm2ILcyYyMpDsDmJCqDscoG0CTQr7KjWiXJ5k2G2lwIUfI+OMFDvk8QYIBnLjEBA8+5n
iCs+/W8rT+kxUWhk7BGtVfkgGbwBqzZYJA4RaaEwgQUGsJAHO954kg9+S+BfeAXGvctNGSdlb05g0dTWJIXkORLJscF3QF5S9Tc1gT6HWFzKiCbRJr2HgYyrX3ljAm2I
2J5S+loXhnzHjm7LpMyNlmdRPIgkffoAyTEEpyWHejMboWUVmVMtK8A9mk3pKTJNQJpUJxl+RIfNOki6VogZ30XPc7K6ltcHTyNhooDlkj5q5DA0/ZFFvZvZcnuA81Sf
miI9362LMLPNZZ9m2lLDRvEzCcJLAM51HsKOUktLISMuiegFVfxlQn6dmFrKobIswEBwuPTrmsXmyWZFoZu3a8qIJtEmvYeBjKtfeWMCbYgmp+CAqR0Q/CcMzLlmizOj
m10kzhbMT5oW0n0QrhPQ7MqIJtEmvYeBjKtfeWMCbYjHyi4l1BMuW9z9RHFERHTDuHQ2dUOeKWtB3BY5yyvE9fYOXjc2w1gU6tZCQaytV0qTP6fBPGYsjJ1Rvh4FCTOH
AcTvF8gwooMKmKArv5m08EXTT7aPrvZJ3euMy42MAF7KiCbRJr2HgYyrX3ljAm2Iyogm0Sa9h4GMq195YwJtiG+DmYjiSRK1MTLi9OAQjpWeYWjzdzwhrNDFY1tx3p28
2/bKtlshAIdjfLyduhFtRqPqArepcrA0lJsScS70YqmX7vm5NZE+NMF42FKUlaSfyogm0Sa9h4GMq195YwJtiNodxBqwmU7O5NMMqs0JYDWtF7e9Suhq6Ph9p+32CUuy
/ArxS/Z166l2bwIqCG9P+53F9MddNVBrC9w18hfiQuXRQpxScJy4aXZr3i2JwQemUaAX7U0hcYZzSVXhat4nBsqIJtEmvYeBjKtfeWMCbYisu1nb8Y1qgIq29LhBJALG
UroyKgW1UTm0M8KPPbmhOEefba1b0fX28iqjSHn31uqOMFDvk8QYIBnLjEBA8+5n84qBee+w44g7SXPBYBuoi1y0yDVNfOwHzVFaczKXlkMCtoIbqs6JW6jRcAATcEwe
ZE5VFl+RXCG9BsyXi2XMh2IhQtAqArJHKkcBoDi2F4TKiCbRJr2HgYyrX3ljAm2IifBsOYHC7REuJipnwHIbY0cKdlCYxfgDXjYXYzltKg/KiCbRJr2HgYyrX3ljAm2I
oPejuWTbTvma9Hj0YVw56Z0bvupPSkv/bkE9dD0OoHI9f1k6fti9G1UtnH/9nXVbh567rvEwS7Ivg6ofhMwRYMqIJtEmvYeBjKtfeWMCbYhaX//m15rZnjMgLugURPKd
yogm0Sa9h4GMq195YwJtiGHaBzt4a8gy31WxvuhMz0HljoJbdqEq+gCaaupRg178Yj+qsCvGSnZQSj3LBUc28/swZgDkTP8lU4XTlB57vs0iSck/qKKk0zZI5JPehSnb
yogm0Sa9h4GMq195YwJtiFiiM/UPb8MeEeONk3N2ya9AmlQnGX5Eh806SLpWiBnfZize2DgwchDa0yOySYRE4XHQOM1gDKFZPNQNGgLTKxrKiCbRJr2HgYyrX3ljAm2I
OS1cgCWoYMf23FjxgsjcOKxq2TGR18WWr8RCJzMH4GXKiCbRJr2HgYyrX3ljAm2IYqtMmuOKAZl/xk6DrOmNGU0myab+Xu+TV+vnXhJKD1vKiCbRJr2HgYyrX3ljAm2I
XPOyDk3IC0mk6GbfpWB41BHq1BIXKbI2En5PqNNNCmhb4NtxVpMbBHY3gZi/tdlcvBXdNnxQ+/ZzgkBbox5sUWROVRZfkVwhvQbMl4tlzIdgdJ/tafo7o4+AbyLiwPuT
yogm0Sa9h4GMq195YwJtiPetSo46JNIh2FMgyDkdWK7/ALDxn0rDA2liWlB5d7+/RQeZghvvbzto2QWmwvOUnd5t7+F0NVq8oxTUtyCQg1aIKAvHqTpI7txakUUmAFch
KW033gHjf4EggCKWz0PfOIVjRAhXPkQhLRHHwEP9y+gxd6VKite2vfN0WCjefC1oneOqIseipfxSSmi4yWoyWiN8bsVPQeppNDPng9UeWXXKiCbRJr2HgYyrX3ljAm2I
G9hykwbwJjywpy92L8RqpMqIJtEmvYeBjKtfeWMCbYicfu3vj+HhdKs/Jsgv7+8tzr0PpUFrGHIEKln0/UyEGwODxd5pDbQ/2WgekQu50rgLdN+aNVl7/5GLHdAaCQtg
yogm0Sa9h4GMq195YwJtiFzzsg5NyAtJpOhm36VgeNQY8/lLiKsZpWyVnQp2VSPGCx49ZDISnGwJi6i6tTbQNqoHj5AKty/a+67172h4B5PKiCbRJr2HgYyrX3ljAm2I
ZE5VFl+RXCG9BsyXi2XMh6UtKrO5gTibPQ4cA1l+uGnKiCbRJr2HgYyrX3ljAm2InRu+6k9KS/9uQT10PQ6gcsqIJtEmvYeBjKtfeWMCbYiSNiP5m6moRQbLFIyOUiSl
rRe3vUroauj4faft9glLsvwK8Uv2deupdm8CKghvT/tAmlQnGX5Eh806SLpWiBnfnifbija+sB8ruJRhqSlUlmrkMDT9kUW9m9lye4DzVJ9AmlQnGX5Eh806SLpWiBnf
Rc9zsrqW1wdPI2GigOWSPtGWBnod7x8eRXeOfivovXPxvSqpKMYOBxXvuIPGZSx0yogm0Sa9h4GMq195YwJtiPetSo46JNIh2FMgyDkdWK6YY/bUEpAjA4jbK13QXXxx
yogm0Sa9h4GMq195YwJtiDF3pUqK17a983RYKN58LWjKiCbRJr2HgYyrX3ljAm2IrLtZ2/GNaoCKtvS4QSQCxlK6MioFtVE5tDPCjz25oThHn22tW9H19vIqo0h599bq
jjBQ75PEGCAZy4xAQPPuZxXFdsdoz94eHkH/bkJZeUdsvMXJG9QLTCD9JQRuufiH/wCw8Z9KwwNpYlpQeXe/v4vv+0sdQ9IRSSIe0MBUl3uz6s4HvoNtgafnSWkCbwbA
UL7dXYAZGv9dwYRlTqGSAgpJzuqvwwHUzVlz1AhLkcCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMDY2rgFm8pL1rvEGx4kX8b7
479J2HnN5bMPBOLJagaePY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMDLWuYfsJ+WYR73orusQu7r
pB3CtMmDYrkQJB13/P20eJmGlDrS73sRBDB+mv4VPHhJ7gpR0SzMUxju0moLEvLFj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwMWoSy11l/ktSZ1vGWfBRaBXEK4yqCIpb44Sg3Q1hjJpj7WoFy6tbRuDSxIbySiAwMzOJ13HROhAr2M7jFs4lSFl/MiX2v4cuhzgzagWuCTu
JMjHbg5sgc5toUk9uRtdVI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAKWhMGB7tD4gfdH++B1seq/dYSAc/nCffYZYg+5YJlq6bXSTOFsxPmhbSfRCuE9Ds
LUbso2j+PvhmQG5CqvWoQGobhh1gAcIdh6vWrgP9nkUgSYyvVtufLF5ns0ScUSSMc4P2kONHgqskGsQRo59xxY+1qBcurW0bg0sSG8kogMC74w4wEBAepOCiQ0nq3dzK
cEARDUwEm7/5ltO3u7bFMckEQGAgtrNvMUgEDrrXfR2PtagXLq1tG4NLEhvJKIDAHj7F3Rz6xogmkhI/T6QCNDF3pUqK17a983RYKN58LWin9T2Tcu84UvKb9X4PiXiI
HM7cPHQ4EsIh7d7NV46xUawSlaHzyQXPdRbBrNwMiRBbNdTc9rMOwrISgUhPI8XqqUDlsHPsOarwjPWDuRNgYltXriayqgNGXhWTfV2b1Y3AQHC49OuaxebJZkWhm7dr
X+DfzUSLQv0FuhERws9LiuAD7oWMY2TKQ0ZTBgMMPYnVOIlio0t8x5Ykqbz54tjhnRu+6k9KS/9uQT10PQ6gcnz7oJxN6ptkxjLYq5F3NsVoYAax8KpR9ordH9YPHB99
cUgCfCi+0d6sOxBl5Kt3Sriqidc9EI3PLbe4vSF+HhTZVy+MNygeHzEN+ZmTFKRRieUi3TEOkftmcjKqfl/tQ6MNZZo3xUZ6XlATG9OwMQPErOx3SCsyLsD01zVjBcdF
EsmxwXdAXlL1NzWBPodYXJ3F9MddNVBrC9w18hfiQuUree6D6YJ4i8cU5ui58tVPY+NlxU8UFuo0Q1jLJxjdKuhrJwalZbFKEc2kxjeFJ5+qHv6lVwapfnwot1m8KMn9
+6H6JzUxjCggCQfNL+Knc+ckAVFMBTXuR8s9QTXd9HLHgUU7MDSqxkjsiwyZgJIROqQqwCFg8Zb1cLnkhSalNjxH74y17RT9IXVPaMmlSMypW517hhVFJrVdRjzBPzRA
er22+NdLhgHNVWPZtxYptB69oMVxh6kgXtfwbcaBcD8xd6VKite2vfN0WCjefC1oIHhErYfIcgTrEjooKVYYTV/F1jNqoLFSlR4tQV6ke7CIBfNNSuZ8AZtomkozMvnU
N7zjCz4Pu2tuZNtfj12k91t/+A0Y4zi+N2GMiH4LDkx+YIkjTcrnYsp44dr9P4nI/TNl9uo8MdNfvgkk5vgaw5x+7e+P4eF0qz8myC/v7y3bJsjEjm0cwM+m6hpVM4os
bjTdLuKg/jPIEDLWxjH+d1y0yDVNfOwHzVFaczKXlkMCtoIbqs6JW6jRcAATcEweScG+Doc6Au3TZfJPcmwCqUcKdlCYxfgDXjYXYzltKg/xMwnCSwDOdR7CjlJLSyEj
eXXSW6XSGLk63+hr6EA4ckvHzBbmplGJxe4xhh4uqJHAQHC49OuaxebJZkWhm7dryogm0Sa9h4GMq195YwJtiJBTt97uAw5szgK2LTcP7O0jMeXwrwUm9EeGeZU9oPTr
/wCw8Z9KwwNpYlpQeXe/v/YOXjc2w1gU6tZCQaytV0rNzOBigsG6OM7sofRpeOomlg2Hj6q8vzdCMoyYBN9xtLo78c2rRor74mCOIT+/uDpiBhriOEqr6cUQpm1V+I+R
TaqJwlWYYjuZjzZqwvlzL3MZs5pjsxCfyQo62I6Td9meYWjzdzwhrNDFY1tx3p282/bKtlshAIdjfLyduhFtRk9/c/uO32XQ7QNsEo8oCovc85vMGbHGSaKK+qwFNOA9
5vF6vnlahjQmkS8vjJJRk13tJwDxg01Z8aqOVt72SgZAmlQnGX5Eh806SLpWiBnfD3rvBhMAyzrkn+ushykaHtGWBnod7x8eRXeOfivovXNibuDieN6/6YLGJ2h3d8yS
E0+AX7xi/f7/1d0Y/VbZDsqIJtEmvYeBjKtfeWMCbYhc87IOTcgLSaToZt+lYHjUZE5VFl+RXCG9BsyXi2XMh8eMe6JRv8OnluiVo8N199DKiCbRJr2HgYyrX3ljAm2I
oPejuWTbTvma9Hj0YVw56fetSo46JNIh2FMgyDkdWK5ozeQugcjwo66MHwd3Txijv6P7IP8UibH3inDccXIgtDQr7KjWiXJ5k2G2lwIUfI+OMFDvk8QYIBnLjEBA8+5n
SEISxe0PsvMzSo5YvmiYCluMwOpps+WrE7F0o4Quyg9ctMg1TXzsB81RWnMyl5ZDAraCG6rOiVuo0XAAE3BMHknBvg6HOgLt02XyT3JsAqlHCnZQmMX4A142F2M5bSoP
8TMJwksAznUewo5SS0shI3l10lul0hi5Ot/oa+hAOHJLx8wW5qZRicXuMYYeLqiRwEBwuPTrmsXmyWZFoZu3a8qIJtEmvYeBjKtfeWMCbYiQU7fe7gMObM4Cti03D+zt
IzHl8K8FJvRHhnmVPaD06/8AsPGfSsMDaWJaUHl3v7/2Dl43NsNYFOrWQkGsrVdKRrb52KDHDJkxcvjiiU2eT+wyl/oMRESf9i9ZGCpHStypW517hhVFJrVdRjzBPzRA
QJpUJxl+RIfNOki6VogZ3w967wYTAMs65J/rrIcpGh7RlgZ6He8fHkV3jn4r6L1zFcV2x2jP3h4eQf9uQll5R0T8slFKZPC8ikwXshEPIdaz6s4HvoNtgafnSWkCbwbA
uRiAYDnR5ziJZmPDOESAhDF3pUqK17a983RYKN58LWggeESth8hyBOsSOigpVhhNWCm+iUaZ6uqqdBpkAxRe2/8AsPGfSsMDaWJaUHl3v7+dG77qT0pL/25BPXQ9DqBy
qekyf2lt4+6QqOLCav8diq7KornOxBT3V7fwqFO9NM2PtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMDpnpEG+56ZBGJEk7psWlm7
uvpR+mDy3ZI9gc7wv9TVc3Hx4N/Dmr9j6r2KunB+nr+PtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAvvWIIJanZhqLlJt2oDeHC
hnKU53E3ivtTsC+q0aEVsZP5SHbn0XXz2m5ZyW0q56HEf9q3D8GeLJeGJc9zAr+pEdbmwgvgU+xW+sO+GBMORo+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwEd8Q/5/qyeLnUDxO6/5m2832wOdy/aGP3iCUWCXKawpj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAO8qLmZlzlhsbVJUFtOz8L
iWwvaOy60QEgXjuWUKhaU2bauLJakm96z9CiboY85v+PtagXLq1tG4NLEhvJKIDAsoOyvigrKC1uDrOpn6cGwCFexk41x8OB3DVXR8zoSto8aNn0aBCHg0mjdFO0QyJD
lE/qCdHjCHqcKuehq+snbL0aYnQI48lQTVrqLLE4tXehoMM0dNozKgv/oqwZ2HBDKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMAmHbIsy7j2vbBolihoIMRX
oiZcykx7AarbX6hjGicXMOcvpR0G1G1q3RMd3JNYoyqPtagXLq1tG4NLEhvJKIDAIRwpy2kiqk7GhTpGZ+SCgwl8QQBgzAEvRMHB9qPR3gKaLLoic6or6VTo3qxeS4Ne
Rh8m4GHFKs3MicUN2tq7CPTfUixbRote9r54PCd/uOB9l4uPSZ4zoH2nlxmUWHNoxz3li9s3n70PJ/5eXZQuw0etQ/ZIAJxfidckmkzBvo5mug67FcZlKFQCsa5NL0lp
Ym7g4njev+mCxidod3fMkt+SYTldFiq0c5L/J5m6qpLjPmBYjq2k4W4KXrkjScX+9JGszkrpz1WXkqq7RTf9LYgo5nqny+DmDItt9IwXS9meZ5mUnCVk0y5mECOiqffh
rt4WMfls2v0IR6labkuEl3va2KL4n0XOmzirwTuukwleOZXMZf0IuGFnbXRAExAGCBa7B85Nx+5Qr3paJG+jT8V6Ik/cazENBOu0wEOFvuNsRj5APzZ1Croi8zbqyWvG
5yQBUUwFNe5Hyz1BNd30cvmigenEvTx+UX/ixClIEtPK2O3l/8k/5f0z1pUai6nnj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
4hvPX91d8/vxuywFQajYcXUZ5IxQXUMQzDMeYYJNWTO751ECO64iAOBsGh43VFR7bHDckEvEh0ctNq3WwhM5vI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwN3rVyZqjz0BAwvpo7dsjj/JAAbaUmE9rscRxUXXirZcaQjDPq334pK5U5VpvcLKE58WnKoqwfnoZNopvZNBn2VfkDB7xohPE+2S7HRhQ80O
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwFFH9EpOysaBSnbWA/eVUhpUwTaEPtHZhcItmdyhIcX2
/8bx5c+/QKklpzqQx/+F6I+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMC44TlwYF54DSmZ7hmUN4re
rWEyM/FszOjf0JXUipSPUJH855IK+ieKAYhq0vZrmXVmo6JXpJxsR/zFvhzFv6z1iGohucOz2F60e4g/fpX4no+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwJ6xVsOuQdDZDY7xXgoKe8CEnt+uw94lQhhzizr/dYmd6+qEacJdQo7pe4GFZUJ3w4+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cIedeMRtJtvs1eGf0/eToKDTNJ49A4ggqoUCwAZvKk1gIlzCxjUxUtpmpnCJs7gZJL6PW0NjRcEiHptH5M5pEoi
aWVuBydEyMzfevhlNU7AZGisHkdOd300SUBo2Kh8Hx0Mr00N5ZD6jmvrY7ldUxNWe28BGs8lN9xKmbAyDdvCcAYsEMP+vfE/kokuMNvqkHCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAytjt5f/JP+X9M9aVGoup54+1qBcurW0bg0sSG8kogMDX0tFLODqgoU5YvLqL1TCO
nSmOYzLAA2TYVR8/LMD6W67KornOxBT3V7fwqFO9NM2PtagXLq1tG4NLEhvJKIDAzN+Lj+ROXQ5LAkTqt3qVxtLAi0t/e6IJrWwN/MjcADSPtagXLq1tG4NLEhvJKIDA
qRj4RwXbXch8rZHvniML+hHw4DFqXSuMUuyrS05CrRePtagXLq1tG4NLEhvJKIDAeG6e6k3u8u8RpFk4tA/VnAIbt40bClc5sB9+IyzWzuKjZzaDkt6wRQkMXmZoGFpm
PXbfNK/bM63pgM2UzllWef9sb4cS9g05MIEEEjulkFLDTOLVbksBK+xKoQ0yGQMqWjLFV852TmX4leCo94HFXIlgLXrPGCyMjwkMshCrm55yaR39CpOEWgNQKG2qMatR
QjdNrpQK0UB38lnR5fZp2EvoGZdZmyIyRMvPttDbReF5BnVMEkgGKA+xnnHLrgesGPABjcaswZQJvHPcULEGzDQr7KjWiXJ5k2G2lwIUfI9Kvzk1Gw8WKJQv9gSfjQ/k
OA9Nsq8s9DTSMjSYDD4hNd+kE25hxX/7mEOCpZYi+aBjch5fTEgBy3cL478npottLonoBVX8ZUJ+nZhayqGyLFzzsg5NyAtJpOhm36VgeNRwbVQT+vz3yvkqCgxEglkR
7ltxsJfopQTr/3U1U6w/x7Pqzge+g22Bp+dJaQJvBsAscZ8v5qb/HX7q+7TE7S20XiMg9e3hpRWm8SaC1KS/sI+1qBcurW0bg0sSG8kogMCpGPhHBdtdyHytke+eIwv6
d36818+gED88v8pgm3trNo+1qBcurW0bg0sSG8kogMB4bp7qTe7y7xGkWTi0D9Wc5knShrhWnRsHMRd1ETTYOZI6xWru8g49Eoe632yObXqoW/As2NPz7srNLv0iCRn8
CknO6q/DAdTNWXPUCEuRwIkTtD4+JQAJdIisJ02TW4xi3gB3q5Qru8586LQ8ZkyOrsqiuc7EFPdXt/CoU700zY+1qBcurW0bg0sSG8kogMDOWiSRndtIejByJbD7idU/
WRvxAPSiVKF3wWD6zs5d/WHyX3w9WDTEk+GlvhSk/cLiKoPLMYe+1N2pnJXmPsp+8PI5dqy5Koh5lEHB55bAKGHaBzt4a8gy31WxvuhMz0FAMlK8z9mDkYfeV7Bi3Zsg
dZzbr1R+bIRlnYaAvHoDhZoiPd+tizCzzWWfZtpSw0ZNJsmm/l7vk1fr514SSg9bqVude4YVRSa1XUY8wT80QPFrVeZsGo6cPeWewF7mRlGRlWaijYz0CrLBFopUaBPr
sAtH8IyqSdxfPbqUOLhy88BAcLj065rF5slmRaGbt2vv1uIBYtGoG4zIeb0/9050/2xvhxL2DTkwgQQSO6WQUulzbubDEjDb0SFepkr+qXNibuDieN6/6YLGJ2h3d8yS
TSbJpv5e75NX6+deEkoPWxLJscF3QF5S9Tc1gT6HWFw5gSQGocpVa+S7ePSWGvk12N48TQBu6FA2iD0tMg6sB2D8Xaiw4ZVJuNhPNIY1Zbaz6s4HvoNtgafnSWkCbwbA
s+rOB76DbYGn50lpAm8GwOXUhor+/mCFuGBpdPrm52dQ0n2RCOKRIssQ2IAol2MbCzaq0dvlsA6RRvE9MXDzEmCy3EpC6x6NnWbv90rW/40bdR89K8QjjRP+TCLT9VHb
BDA3WoLuE+nc+UU4bIq2eSjB45bpHUM4lW9Yc29yYoEePsXdHPrGiCaSEj9PpAI0Xru4OAGz3Rt0yj4G/kXNIwpJzuqvwwHUzVlz1AhLkcCJE7Q+PiUACXSIrCdNk1uM
WzXU3PazDsKyEoFITyPF6lKGG0JF9gH2+6r3RtN/te2KhiY87QWvZ7rOnhbq8sNywEBwuPTrmsXmyWZFoZu3ay5rcjXBITqiOzldN+flmRvkpzOzrG7dcVYb5TZMXped
XPOyDk3IC0mk6GbfpWB41HBtVBP6/PfK+SoKDESCWRHuW3Gwl+ilBOv/dTVTrD/Hs+rOB76DbYGn50lpAm8GwLkYgGA50ec4iWZjwzhEgIQxd6VKite2vfN0WCjefC1o
CeJUlNwRF6eJh7C7uU01R9w4MB6ZoE5Ic0BmC/dHkHrxvSqpKMYOBxXvuIPGZSx0miI9362LMLPNZZ9m2lLDRvOKgXnvsOOIO0lzwWAbqItYojP1D2/DHhHjjZNzdsmv
030fEYbTGltZy34BDLVR4gD5HxARTe3ntUngb6ffQATynTFmY3pQ1PkTuuPeJCISytjt5f/JP+X9M9aVGoup54+1qBcurW0bg0sSG8kogMAqIMH4mgFS8m5cr+mr5RN3
oyGEfms+tqtFOzDWJyZdKI+1qBcurW0bg0sSG8kogMDzBc0tCsKRFUJDp9JUP3rPviPBUfMABYZu2PJ9sFxgbEP81Ha7QVdcjtviNOjbo1QLNqrR2+WwDpFG8T0xcPMS
YLLcSkLrHo2dZu/3Stb/jZz3Eyy6WafSKVRbno14G1njr+j5usfLNOV6Urq1/jyAMXelSorXtr3zdFgo3nwtaEAyUrzP2YORh95XsGLdmyDJO8uuSFifETujQUajQjuj
Ym7g4njev+mCxidod3fMknS+/hyH8aLnjf2A161DSDuPtagXLq1tG4NLEhvJKIDAdYgqyj0nFoi/OdO2gQsJSJaRwhohdYh/6VR3ZPom5p2PtagXLq1tG4NLEhvJKIDA
PFV72em/UtNMcRGCClOi/Sy4GZeoKjoyDGRspFPolKI3P5ElahsOCnM8PE6X+xWOWKIz9Q9vwx4R442Tc3bJr+PxdrKWukKprGVrusN6t8cxd6VKite2vfN0WCjefC1o
CeJUlNwRF6eJh7C7uU01RyYa+CkclJxEJs3yvJ1MFwLxvSqpKMYOBxXvuIPGZSx0E0+AX7xi/f7/1d0Y/VbZDhLJscF3QF5S9Tc1gT6HWFxVTWLC9WyYvZGCtr+g8wNY
MrR9m/PkGyDd9ht2zwvZN8saR6u/UFMOHQkX4PeuEhvbCNwKZQf6ab0E2f1jdinQpHk4pyaNQbN5K4yY6gmiNFs11Nz2sw7CshKBSE8jxeroMz8cCm0njmXnMMBWcNvL
yy8FTmQEkQyDytWnLZwM3LPqzge+g22Bp+dJaQJvBsBQNdK7/FgOXJlVBvWYhKdcj7WoFy6tbRuDSxIbySiAwE7ITT+IFtCIJc6nr7kc2dxrGa+zlLW4snUM1QZu2Sjb
j7WoFy6tbRuDSxIbySiAwLKDsr4oKygtbg6zqZ+nBsBaQDM4kwRzq51LjjXYGgU9SAIjJZ7+CPk7PZ9GYvFtEmHaBzt4a8gy31WxvuhMz0EvQw+s0QUAizwSRvI7/stA
+tBLqa3rGvI7blMlM+rvAMcp8UR1ywOtnbZ2c0OxBvcAjPNiQ97jOo7wV4PS92HT8wyh1OCLzUJ9Fwbsk410tZElii1cozzcPOcPtUciWKhk8zLP3nMUB3EsT9hoPdmH
1R9fgKs3gvvsG3p00hJwFI+1qBcurW0bg0sSG8kogMAUKCn2/qSdR0lHSaOSgLLl46NDeAoOrWvNGxDF+2YLejZ330xoUcj7QJN7ORy7OxfK2O3l/8k/5f0z1pUai6nn
j7WoFy6tbRuDSxIbySiAwABFMY50SBmF86+73PURyYFvsQepjPswsjPN/UUcpF2FZpDIIg0rnfUm5tfmJkQM2touYnTj+L6K9vdV/hxmK/qDsvK+/Jt0twIy5NnLF+VG
KMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwD+WlZhTnZXN7JuIJFDHwQl4q+vwI9AC7T/AASGC6rJF
ytjt5f/JP+X9M9aVGoup54+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwDAxFCqvcjleHpxggUcQ2HjKYU8u1ZH57YqlNlPfhyNC
rlkb/I58jfuPl5foNt3WsXCiBjYjsqg/i3QdygNer1tzg/aQ40eCqyQaxBGjn3HFj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
Yzo7S+/XGUYuj9JQn3nuYy9TC+PVR7Ebe+C8+bq23EGPtagXLq1tG4NLEhvJKIDAHj7F3Rz6xogmkhI/T6QCNP7K1+bpJmsDvZZ0Syxjnsd63xvi6GlEUJknxEfSAgvt
CknO6q/DAdTNWXPUCEuRwI+1qBcurW0bg0sSG8kogMBKYTRDgMVBJHeNlvVYNYl90cjbXh1VGdHq3LvVUgtsXWL0RBrXRNyC9VH6oA+bratFzWzUaKBvUZA48U5VUZ99
vRpidAjjyVBNWuossTi1d6GgwzR02jMqC/+irBnYcEMoweOW6R1DOJVvWHNvcmKBj7WoFy6tbRuDSxIbySiAwCYdsizLuPa9sGiWKGggxFeiJlzKTHsBqttfqGMaJxcw
5y+lHQbUbWrdEx3ck1ijKo+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKDCXxBAGDMAS9EwcH2o9HeAvnERbYXKjtM4YUqKLi7qzRq64LFl66SFIDMbOTJ+7RW
gz6NJ3qq7K+KvamdoL7rNMJd4yRouVe82Gpvhgn7crLcecbOgewXwS2ciW96c1fE5yQBUUwFNe5Hyz1BNd30clSexGWuanzzxHEOAuPtBmucfu3vj+HhdKs/Jsgv7+8t
AkAPLKUdYyX9AjE73sb8/biihoSvwFmKMImRLicwVDe3xg0qClt3JmXafxRI+a8kRVVjJBx66Bd8hHBAxMSwsGOj8BZCOR9K1ZR+51aVLJN6bpeBly/RF0SO1jOHa1vw
/3ZeYJ98TVOKOdJnkGGCk8aWs7e0lxC/yyqWVB4y26/KxuSlzMDsk1OHw08yTJT2bpNAGyEI2ULqKnSHZ1omAIEh9Ur6mtauNbdP1NuqwnXioFpBX3YvmfTdMzYpQveg
i2jjPF9b9F/yY+yGZnP9r4+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0Zn2Q7srVwq0PBnosfMIkAUGiMRI/R7wWkNhxsPVfraeQzPrtrFfSIZRyiMCKoShP
i2jjPF9b9F/yY+yGZnP9r4+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0hsPpradLEdyhiuLcyOKNrDx12youXHKa4L27mzUTHtJJTaM64u87kwd0hyizCU+A
tW3ZQRBajtEWRgMCpSVpUUAF7ZqSxUOfUbnENkLLUO3o8ap8VAgT7nxJFqLtMF3wYrobmFH7J1+BahSWHiKg4o0YPDIBb0AcyzBiq894jre25DK4207nQrojviTuW4mP
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAdC0TjMwbz2VY2j+o5HP+fUQwAdoBOC8wBkU+1fezGitY6FFv8WBzJxjiKupOkLycztgnQ67XzKqKKV68/U5kB
fNgrzi/S8fEZDhomekoRUo+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAjjBQ75PEGCAZy4xAQPPuZ5GfrgBXc2YhK+C/rowi0q5vjT2ok9SJIzVgvmWfNB37
i/ySMCvL3lAYbSEiIZOiIO/W4gFi0agbjMh5vT/3TnRxMZX06I72LO1Izrkg9auVUklbicqAxfG6sco73kepbhC2e0e9QmUnyRsgeikEdQ9ABe2aksVDn1G5xDZCy1Dt
pndvazvkC2jASHlAB/I6mSlLbdL6LBDLNUwX6bJrqQmf9Tx8GXuEJtWHN3BDbOpCVU1iwvVsmL2Rgra/oPMDWHAZXh+V6gagR63WfXPbaSpx1Eud48tj0y4RPx8ae8Uw
5Ov6Ep50vcPUTr+qGMVnMNPQNDU/3oZawaMDNnnOgAYQXo3+wTyO+HudCMiaPfi08zjY7+s/mRss6w2jg+DmEExAUUdAwmH5KNoMfp98lh2f8IRiovqXqA9Ixp/APU7u
OTvqvI7Ihg8NR/E+GFxcoo35L2C7eXjXtnh4N0eGmKnAsejAtKlZTUfRhc79XdOVTZKSFnzf7wygCmqxHDREIDoFszDF8upN3iArgsZe3JtwTsF/Uet4hAMr/vcMDsDq
Iq10aZRpV8R7us6y0zouVNMAb/ZmIp+g9tXlp6kmkNKw0l/dzgJ5Cfaei1uMxYkAKdRqe+oJe0bnf542dn5r6Ds5O/J5GjsVYBUPfOKiCgLEIF4GmgdSMUZkh+UVQQ4F
IXQkLYgFVVq4adXr0zhVGB5FLr0IMTWw4utSDQHcp7xJld1HA3ixoQP+zzXD+t1MTG9py7PsR6VwxaRrXjRRjskKh+D3K3YJSN8zpkS7pT4+Tue5sSXeu74wJpbMw/c3
1d6JlEeD2G6sNbXIQ5zFFfPRxMrqNk49+5Bhg7DXK/CPMb+MXOr4+fUdlu5UTtedZ3xJmfiVofyKcdiUbZ+wU8ZwPcu2fWGvsqh72eP5lyagL4TkOzLS45wNti6nXcKe
SNQ+ij3SacI8MlyLHNrrimI/t9wc53hL0oqQmhqD1DYZKcCI0koqMJIJhlgcm6L2nRu+6k9KS/9uQT10PQ6gcqnpMn9pbePukKjiwmr/HYquyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA5H+Ans3CGAHUPj9kzKm0VMNfnEJE5w7b3ycaNYkcNlePtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAqr7yffXqtJLzZ2o9D9uH/gVxzOXK/717jUciNWQNQrwZ4h0FZ2xER61arDJWTXKs
PX5I9s9Dm079D3bKcWfx5BUXivM1n771Hfkg13AwwodDYBrbonSZRXZm1MiGEVzMMf1Sh9MojdpIr1ITEWLzULS98OUCEHZYANZ8tliD7MwEE6RXfpBsxnuenZkvPqTu
fdKgoISTa6Uwgy/MA/XCzMrY7eX/yT/l/TPWlRqLqeePtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCxTCRvyHw/qIYM24uwdmVq
j7WoFy6tbRuDSxIbySiAwCQ3iDsa26VCbi7qBViwuHdqd3pkYpqPPwYmNt+UmcJLYDoB9k9rh5Mdk9Mqg1VvOI+1qBcurW0bg0sSG8kogMDn+fXuG+gdwubako4MCjwh
ApOYzFAD6+QkvBhI+gBLWS8z6ZKuNYchV+GCWpt2+pcvM+mSrjWHIVfhglqbdvqX4o7HpnvpjVTcEyfQXJ4ifDLstgycJjKx2eTA+Jris3fB0hcTXmdGpPGzksxappjF
LzPpkq41hyFX4YJam3b6ly8z6ZKuNYchV+GCWpt2+pfcZy76kuiEeRv63JQWy8iAj7WoFy6tbRuDSxIbySiAwB3iBscbxtpVTang4aPXCEjUlm+VlETJi4RqX4r+wqfF
j7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cJdPC2/E6r6xENby/8VoBQD9Gt30COWkYM8T/Dg5IKBM/bxciNBDLtlNVcarSyAxI9VXPDQXzNE5gHld1Pl/Hcr
qVude4YVRSa1XUY8wT80QMH9M9LkPYEX5+lm5cjtOyLKiCbRJr2HgYyrX3ljAm2IwDD1ZvgMERTUCrVmf8kQCr4UJ46+rd/lWRFg7zB2oukB9+dOj3WWisinHOuvTsYo
/ArxS/Z166l2bwIqCG9P+7a8FJzqwNUx2xPq1l4QEac7JQca+gE7iqg9kjbO9ja+5SQzn3scf6MVONfjzxq+c2HaBzt4a8gy31WxvuhMz0GiUBGojsYltK0rsP34Mbh1
4J6JS7+T/oJTjj8oLvRrWvYOXjc2w1gU6tZCQaytV0qKayykNAYT5yvrj4kxFQ3aWstj+K+E2UODW15yXBS5K7fR3CF3R+ZkqICUHy7gHk776jB0XKTasgRWOT9xOXA1
/xKVZtreaQx/tCmlzC6KXR7ORmfm281/QtLu65OYUgv+Hvsh9YmjKUfvUiN3aUnunRu+6k9KS/9uQT10PQ6gcp0bvupPSkv/bkE9dD0OoHLHgUU7MDSqxkjsiwyZgJIR
yogm0Sa9h4GMq195YwJtiMv27KwTyTqMg3d9cHEO83FYdOqXATaHv/u5ice2ZP8NNCvsqNaJcnmTYbaXAhR8jxKGCCs8v9ykxoyEzgTOIAtuPt2lzp30bcpdptza/rZT
DAJVEqiG7ZjYaoAe3NPboZ5haPN3PCGs0MVjW3Henbzb9sq2WyEAh2N8vJ26EW1GusM+xrjmFXFMEtZOlBokltc+zZqcVimC41fLIWZFBkn/ALDxn0rDA2liWlB5d7+/
+WgO2/xOkUC/oTHKljiwG8qIJtEmvYeBjKtfeWMCbYhBNV6kO7Gtj6OJti0TAY6GwEBwuPTrmsXmyWZFoZu3a+/W4gFi0agbjMh5vT/3TnR4Iz2LF9Uzk8Rc4ULWc0H/
yebSFJo7ZOCGQP/SCCa60PetSo46JNIh2FMgyDkdWK73rUqOOiTSIdhTIMg5HViupFGWZYx13hx5h/riBH0tgo8xv4xc6vj59R2W7lRO153Ew397IJG3SzIt3fhnXCMo
xa8cOJHTF37f5Eq3NkTiE5OhWaO8oeVjlF7c0bS7Cisg/z1fHLO3jnrSplZ+n/YByogm0Sa9h4GMq195YwJtiPnHB86ilx7uzKslbgO2HP70d7un807p5FqkeIFcn3b/
mHSJesLcxZ5Sg/2/21vqbxs9cfr8Ks0YuRO2YF4SfKdibuDieN6/6YLGJ2h3d8yS84qBee+w44g7SXPBYBuoi13tJwDxg01Z8aqOVt72Sgaex+qGqEmxBXTeDvDoM9Jq
J/4quENb86UHz1iWRxy0uYvv+0sdQ9IRSSIe0MBUl3uz6s4HvoNtgafnSWkCbwbAUDXSu/xYDlyZVQb1mISnXI+1qBcurW0bg0sSG8kogMBOyE0/iBbQiCXOp6+5HNnc
Gpzvs5qtfSbEwb22YuW86Y+1qBcurW0bg0sSG8kogMCyg7K+KCsoLW4Os6mfpwbAWkAzOJMEc6udS4412BoFPZL7B3skzyV6V0aQohkOYQQFSxRDXTjMxYfvHxTkBbHm
qwV22OYXK1KPG0srI7iAeF3tJwDxg01Z8aqOVt72Sgb5kc1W+4LxiV8iqGxDjKuaZn2Q7srVwq0PBnosfMIkAfvUGyGATFv8LxglYIikBvjXBkg/IielxugDTAnqKu5D
NCvsqNaJcnmTYbaXAhR8jxKGCCs8v9ykxoyEzgTOIAtuPt2lzp30bcpdptza/rZTDAJVEqiG7ZjYaoAe3NPboZ5haPN3PCGs0MVjW3Henbzb9sq2WyEAh2N8vJ26EW1G
usM+xrjmFXFMEtZOlBokls3RIA/Iw2Y6LiEdLxtaxL//ALDxn0rDA2liWlB5d7+/+WgO2/xOkUC/oTHKljiwG8qIJtEmvYeBjKtfeWMCbYhBNV6kO7Gtj6OJti0TAY6G
wEBwuPTrmsXmyWZFoZu3a+/W4gFi0agbjMh5vT/3TnR4Iz2LF9Uzk8Rc4ULWc0H//BmrN0le+THSJKBTVcMDKfetSo46JNIh2FMgyDkdWK73rUqOOiTSIdhTIMg5HViu
5Gs3/syKCyw+0yaG8sUufgawkAc73niSD35L4F94BcZUTxkESPYGFVHm8LE5GcCyMHlWETWiZ6FsHqSHNpQ2ZKlbnXuGFUUmtV1GPME/NEDEw397IJG3SzIt3fhnXCMo
S5ekHqOxbhFvOfXunYdzIBeiWDyTz3OZyScvGHP5Upg0K+yo1olyeZNhtpcCFHyPjjBQ75PEGCAZy4xAQPPuZ5RDK4Hdxyv2J1Z47mUlf0lmdfEC2wkAqlNTPhq7QV4b
s+rOB76DbYGn50lpAm8GwPd3qRPNSnPj21Kc7ssCHJs4QaZAOvsVW+kk/dOYU/lfpSsfFoknFbuHwrD40M7rTzF3pUqK17a983RYKN58LWgQXo3+wTyO+HudCMiaPfi0
o2wYMWqlNAyvw8SMoS9+8lsZdQAtdPKJrmJ1Jtq/1+8U4ThECmfSFye2QBoBHK2x2wjcCmUH+mm9BNn9Y3Yp0KR5OKcmjUGzeSuMmOoJojRbNdTc9rMOwrISgUhPI8Xq
JSZw+/a3rIaBDZT6+VFExGN0f9Z64h7nzPZdeNgOl/ZsHMf5+LkmoYQy3ESaD5vxzGr5PmJoM5b2hJtkysEKYmZ9kO7K1cKtDwZ6LHzCJAF6/pq+5iPQ0d8JeiQf7qlk
iVB7xAjAnOYR2Q4P3cuOtHgjPYsX1TOTxFzhQtZzQf9EDPMq9S9hqC6fdj11HJ45Y3IeX0xIAct3C+O/J6aLbS6J6AVV/GVCfp2YWsqhsixc87IOTcgLSaToZt+lYHjU
mHSJesLcxZ5Sg/2/21vqb71322WDa4Ejnu3n4a77/69ibuDieN6/6YLGJ2h3d8ySbRJhH8GSN1DOAUhQGJLVcNC9tCyehhJfVmMkd0QKezCPtagXLq1tG4NLEhvJKIDA
E+gp4cruzzYUsa942lLnv2T5ifwr2JGmZX7TD+f7+1OPtagXLq1tG4NLEhvJKIDASmE0Q4DFQSR3jZb1WDWJfYRe7bd8v7QxJK6Ben040NDoBcfeNIqDDehFWAru6oh8
XKp3NW+FyoHFwAzwfIj1C63lcYcYHQKhvqwuxFZXwZOjoEkZ/V9OyJ6i7IcqBDWVeFuq2js7P6XuCmcZ4BIJ0habKEkXQjvbuWm2HZSnjlj94MuQ1dME7wmxsSfyvcOL
WKIz9Q9vwx4R442Tc3bJrwPjzJB4N2HuBOfxOqogUpRsW2gLNwlOcdMVHe6WLT4Ms+rOB76DbYGn50lpAm8GwEJnYCVrQExOyfuPPy+FWuo4QaZAOvsVW+kk/dOYU/lf
pSsfFoknFbuHwrD40M7rT2HaBzt4a8gy31WxvuhMz0G6wz7GuOYVcUwS1k6UGiSW6dpWFkL31L3iGK9X8U4pxp0bvupPSkv/bkE9dD0OoHKgL4TkOzLS45wNti6nXcKe
SNQ+ij3SacI8MlyLHNrritPz/Tr9T3jLT+XNErsOA6+1GwaxsOd8UYYLe3DW79MxIKkkM1KLIodm0PJ3s1iX867eFjH5bNr9CEepWm5LhJdvwhIQZSe4GJF/zkXNQngH
Vkeka3/bhjRK9oH3M6n1yBXrALABzc6F8H0OqBbgN6EWSA0dyNIYEF/Z4lWPIlR+fSDf8QFUQfSHhQ4hdG3SXpoiPd+tizCzzWWfZtpSw0ZNJsmm/l7vk1fr514SSg9b
qVude4YVRSa1XUY8wT80QILEJGehoxOgc/jvDSGtKcbxzkuQ7bX8s6MCOalk+yk/f1XmWeKMuMWfg7yuQhFDZGGL0ViS/C2p2MQ/nlIRTFKBT4XmyZHQ8Nqvvc6FiOVu
j7WoFy6tbRuDSxIbySiAwB3iBscbxtpVTang4aPXCEjM3jpm/6P/sy+o2Cq/2MT0j7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cJdPC2/E6r6xENby/8VoBQD
9Gt30COWkYM8T/Dg5IKBM/bxciNBDLtlNVcarSyAxI9VXPDQXzNE5gHld1Pl/HcrqVude4YVRSa1XUY8wT80QNf2O6ozYYyVDhDHTIfJqZRx8kqPXsPxv5UQUi47v0ub
F6JYPJPPc5nJJy8Yc/lSmIlgLXrPGCyMjwkMshCrm54QXo3+wTyO+HudCMiaPfi0zVExJ1TC1M+08OxNS7AoaXSQC5vfaCZW1iFACuwqc5g48ElFOZCcsHuLMpZoMpWR
yogm0Sa9h4GMq195YwJtiLfR3CF3R+ZkqICUHy7gHk7AQHC49OuaxebJZkWhm7drCW7CEm+W+X5QSwK8WKOd9lrsE//uHs5tdxeW7tkkeDQIFrsHzk3H7lCvelokb6NP
N5q+XhL9gmVuQmR+a/eeXU0myab+Xu+TV+vnXhJKD1td7ScA8YNNWfGqjlbe9koGx9C77f3yweNSNu/ujGtIOVNj0U7Ag53DaWd8A43vAOdyN5/ptDOxMlafqpGYeDyW
lY43zj+bVwoE5+J7qXikUzSELJjugMpV16HSYYMRLT4AwobkklV8WqLfE9vrAfDMCW7CEm+W+X5QSwK8WKOd9ltGhzTrwZ7pGMHHij/W608IFrsHzk3H7lCvelokb6NP
wC6SXHYPKxRIOeQ8ntsvsq7eFjH5bNr9CEepWm5LhJcOa2oc9Vv0JZ5YgTfDtzv2zHdy9aCYTIGId1IytlH3zTXgq6giQ3e1GlC6olSA1zwVxXbHaM/eHh5B/25CWXlH
I2sgtjyFFtHxAO+XDfKnL3OD9pDjR4KrJBrEEaOfccWPtagXLq1tG4NLEhvJKIDAPaJkxt8gguADBBIM1/xt/I24fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDA
nley/lFqKqRcuafeEUotolHvqV+8S1PU+hW+2moaK03S87gVulpRF5i1wznnkDTksPsJwEOb6Ay6O71habeZAeSRSh/U1s4ejwV1imWTwknT8/06/U94y0/lzRK7DgOv
0qQhC8K13o++Agid6lT2fxzgojoXxykAm/rAluvGF9JdM2+HT7R0ZEwnZe5fRbBh/ArxS/Z166l2bwIqCG9P+5RDK4Hdxyv2J1Z47mUlf0mOZ6TxDBPE0ZVyfSpIGD8U
AcTvF8gwooMKmKArv5m08NcFPjDJeg9/EphFXYqEyjJQhUicpqC1Ojhi8EhfJt3loesYma0BlnQgjoQtW0MlY9v2yrZbIQCHY3y8nboRbUYezkZn5tvNf0LS7uuTmFIL
yhHmAUzeq7gFVrdxrV5foPetSo46JNIh2FMgyDkdWK6kUZZljHXeHHmH+uIEfS2CjzG/jFzq+Pn1HZbuVE7XncTDf3sgkbdLMi3d+GdcIyjFrxw4kdMXft/kSrc2ROIT
k6FZo7yh5WOUXtzRtLsKKyD/PV8cs7eOetKmVn6f9gHKiCbRJr2HgYyrX3ljAm2I+ccHzqKXHu7MqyVuA7Yc/vR3u6fzTunkWqR4gVyfdv+YdIl6wtzFnlKD/b/bW+pv
Gz1x+vwqzRi5E7ZgXhJ8p2Ju4OJ43r/pgsYnaHd3zJLzioF577DjiDtJc8FgG6iLXe0nAPGDTVnxqo5W3vZKBp7H6oaoSbEFdN4O8Ogz0mqAUYXStM2tT4prJQXrEpT3
i+/7Sx1D0hFJIh7QwFSXe7Pqzge+g22Bp+dJaQJvBsBQNdK7/FgOXJlVBvWYhKdcj7WoFy6tbRuDSxIbySiAwE7ITT+IFtCIJc6nr7kc2dz8TbRtPmoqNsbkDEhQ48P5
j7WoFy6tbRuDSxIbySiAwLKDsr4oKygtbg6zqZ+nBsBaQDM4kwRzq51LjjXYGgU9kvsHeyTPJXpXRpCiGQ5hBAVLFENdOMzFh+8fFOQFsearBXbY5hcrUo8bSysjuIB4
Xe0nAPGDTVnxqo5W3vZKBr35+sQOliLqSnsGVSmHtLpmfZDuytXCrQ8Geix8wiQBQsf8Tt9f8ILE+0NqfEU5tTF3pUqK17a983RYKN58LWiiUBGojsYltK0rsP34Mbh1
43KX9B0QocURPgABaybQov8AsPGfSsMDaWJaUHl3v78gZOe6WLLAzMFob2TIRpgwyogm0Sa9h4GMq195YwJtiEE1XqQ7sa2Po4m2LRMBjoZbNdTc9rMOwrISgUhPI8Xq
3RJIihne0T6MOJkYjB75BE78eDnSv86hBGZw2WmJAvHxvSqpKMYOBxXvuIPGZSx0miI9362LMLPNZZ9m2lLDRvOKgXnvsOOIO0lzwWAbqItYojP1D2/DHhHjjZNzdsmv
jrqFRiOgjHW/b6TIYR6fhiVhuqsQK4vU3ouU8jHcqwu6YoHVpJD5cdqdMj91W7A1AY+CGuUsJL5ZJNMN0OmIEyNkuNPFdLIzLzrJMvhkCODHhCnkOJ79KQNeCYx0oGqX
gsQkZ6GjE6Bz+O8NIa0pxnUt6G9cqRAMZtFhidm2dM1/VeZZ4oy4xZ+DvK5CEUNkxKzsd0grMi7A9Nc1YwXHRTQr7KjWiXJ5k2G2lwIUfI9Kvzk1Gw8WKJQv9gSfjQ/k
4yxyLl/l06g0ixpRTiLUbIX8SybcU5HJSTFoHEdzCv3bCNwKZQf6ab0E2f1jdinQR2NvtQW7nCs4O8nPs6/X5ApJzuqvwwHUzVlz1AhLkcCJE7Q+PiUACXSIrCdNk1uM
0D+wCxhqg9czSSwfv+rtha7KornOxBT3V7fwqFO9NM2JE7Q+PiUACXSIrCdNk1uMWzXU3PazDsKyEoFITyPF6selXZnExWdwvwV3H58cn4rod10bYhGbEMqy9+Rj0rea
BNr+7vfHKVmEVC64ZZHLJfc4Xq3bd7Ro4ntzWX+ni8D69juXf6pTzPq3QJYk7+/NL/1JP9Bgl7e0ww9T6PX1zpe8uQP2gtRkkHsWTbo3KjQnHAjKRVwWFV6n1LKpJsf5
NAn9n0QozOeceqVUl4q0WzQr7KjWiXJ5k2G2lwIUfI9Kvzk1Gw8WKJQv9gSfjQ/k4yxyLl/l06g0ixpRTiLUbCHWOAsKzKr1xR+BfCgpbyp6kwZo/AEqx+IEuuWqYrkW
Wstj+K+E2UODW15yXBS5K5cDOw+i8WL5otBI+g1ZKO2jwL09XL7cfeFwGPxPF0wU/ArxS/Z166l2bwIqCG9P+6kEHnz9Lgc19SeliZ20ix2mQyweYeCc/jPle8PgOrvw
YhEY4vJv8+REudGsSIg7bkmV3UcDeLGhA/7PNcP63UwBc04q/vw1SfhT8XrhSr+qNCvsqNaJcnmTYbaXAhR8j44wUO+TxBggGcuMQEDz7meUQyuB3ccr9idWeO5lJX9J
Te0IJyilCM8fKF+tkGQegbPqzge+g22Bp+dJaQJvBsCQsuoNBMFG2d3S+MfcyTVONCvsqNaJcnmTYbaXAhR8j44wUO+TxBggGcuMQEDz7meUQyuB3ccr9idWeO5lJX9J
d8NwmncIGd+Jsa5PGV3rD7Pqzge+g22Bp+dJaQJvBsCz6s4HvoNtgafnSWkCbwbA5dSGiv7+YIW4YGl0+ubnZ1DSfZEI4pEiyxDYgCiXYxvH28yHMEMgSsG88kWXuR01
W0aHNOvBnukYwceKP9brT2TzMs/ecxQHcSxP2Gg92YfVH1+AqzeC++wbenTSEnAULzPpkq41hyFX4YJam3b6ly8z6ZKuNYchV+GCWpt2+pfijseme+mNVNwTJ9BcniJ8
DrW7Q9cXivF1S2ztuD21udHuJUWojegLJYZTo0S8Vq0vM+mSrjWHIVfhglqbdvqXLzPpkq41hyFX4YJam3b6l20lq5kAyQ0xAas7/v/+wUGPtagXLq1tG4NLEhvJKIDA
TshNP4gW0IglzqevuRzZ3I2I+ljkURg4KU+4yr5hn/uPtagXLq1tG4NLEhvJKIDAsoOyvigrKC1uDrOpn6cGwFpAMziTBHOrnUuONdgaBT2S+wd7JM8leldGkKIZDmEE
BUsUQ104zMWH7x8U5AWx5rTc1Zibcm3rpMQ3qozceg+pW517hhVFJrVdRjzBPzRAaigxU9eIpVHiyRuWL4T9cjY2Jfa6PAzwpHF9E2VAsGzWQ3iAxAtKNwt6eUqsh05X
53WdMkHNQXMYTULVBubPQo6FBYfQd31o6QKKsLwIv5I7o09fGceTwIKtOhDsC8wyB+bvUtxduLXRPeNUz/UXYKz+yqLaCeRgd6JQx5yLXfwNhoFiy8FETVBKGSCFGENI
mHSJesLcxZ5Sg/2/21vqbxs9cfr8Ks0YuRO2YF4SfKdibuDieN6/6YLGJ2h3d8yS84qBee+w44g7SXPBYBuoi13tJwDxg01Z8aqOVt72SgZujBhD4J7GJGvif0Q4GiG1
9yNr9aAOh5P+jdDvwvgUQeKHpL2oL4rGZiYfr5tF4fzZaZrwbIi+QDyhg0rgSwRCWKIz9Q9vwx4R442Tc3bJr57H6oaoSbEFdN4O8Ogz0mrf1CpULTX3fmdUlE5cjFl6
R59trVvR9fbyKqNIeffW6vHwzokwm0CiwYmgDmJf+Uze2DfolkiNM3wPtVD1H9WyKI6em2VK8rTntfzBS1o5AHoU0l8EMBvDotqDdivd7hv76jB0XKTasgRWOT9xOXA1
/xKVZtreaQx/tCmlzC6KXR7ORmfm281/QtLu65OYUgsJ+78nEovGfc0K76j7nZp9nRu+6k9KS/9uQT10PQ6gcp0bvupPSkv/bkE9dD0OoHKgL4TkOzLS45wNti6nXcKe
WubRLXXlI4o84GsiPUWNIwawkAc73niSD35L4F94BcbZD2FO+FoKcvGDMhkd2TN6iWAtes8YLIyPCQyyEKubnqJQEaiOxiW0rSuw/fgxuHU/xmguvoycroVpzJ/bMQeS
nRu+6k9KS/9uQT10PQ6gciHslC2Po41lXaPiVPA6SxePtagXLq1tG4NLEhvJKIDASIvAUH/aoTwo2zl76xPodcD4zyACqu636b6Q4IiDCXOPtagXLq1tG4NLEhvJKIDA
zM4nXcdE6ECvYzuMWziVIYj46BF3WFNaMgKSP+OdPdzjLHIuX+XTqDSLGlFOItRsfQtX4z7LadISOGStXi14oY24fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDA
MsiFxuxcDKaOVW+7gHICScrY7eX/yT/l/TPWlRqLqeePtagXLq1tG4NLEhvJKIDAAEUxjnRIGYXzr7vc9RHJgTonwrQ8MN50dQx5gr0YrOI3ht7koiV6KGOm6aUgZUyY
CnA/nEt+4KSJzFcg6GnF4x+xVCPDutQByTTdI0FEZIZYojP1D2/DHhHjjZNzdsmvjrqFRiOgjHW/b6TIYR6fhiVhuqsQK4vU3ouU8jHcqwu6YoHVpJD5cdqdMj91W7A1
AY+CGuUsJL5ZJNMN0OmIEyNkuNPFdLIzLzrJMvhkCOACK6ytcEe46efUzOXePb8t4QDzBd/ICW6fWRR4SCYqC7rDPsa45hVxTBLWTpQaJJZPaKArBgNAXQ0mqY4v27zI
nRu+6k9KS/9uQT10PQ6gclSexGWuanzzxHEOAuPtBmtbNdTc9rMOwrISgUhPI8XqWG11Ka4YyoFbMdW8A8CWpVYi4eqQVITv9/7jF+mhJQ8IkYU2nPEFlBoHDPHvToaS
Lo4u2GmWbL1Oh9j8CBF3Lpx+7e+P4eF0qz8myC/v7y3dEkiKGd7RPow4mRiMHvkE26TmnhtP6aV29Xw/3kRGCPEzCcJLAM51HsKOUktLISMeDaN7NxcJ26ZsCMFePVO9
WubRLXXlI4o84GsiPUWNIxzgojoXxykAm/rAluvGF9K1pNbh1gWFwUS0sqiDECh6rRe3vUroauj4faft9glLsvwK8Uv2deupdm8CKghvT/sD48yQeDdh7gTn8TqqIFKU
8huaYpjkK7ZJqWud3WwFmovv+0sdQ9IRSSIe0MBUl3uL7/tLHUPSEUkiHtDAVJd7s+rOB76DbYGn50lpAm8GwNcFPjDJeg9/EphFXYqEyjI4QaZAOvsVW+kk/dOYU/lf
z3MG/OAnWXwcX2tKs8CBg48xv4xc6vj59R2W7lRO152CxCRnoaMToHP47w0hrSnG3sJ9H0yyl4p8YBWpNCiQZmGL0ViS/C2p2MQ/nlIRTFKBT4XmyZHQ8Nqvvc6FiOVu
j7WoFy6tbRuDSxIbySiAwB3iBscbxtpVTang4aPXCEh8x1xJhrAjipQTLCZxJkoJj7WoFy6tbRuDSxIbySiAwC+9YgglqdmGouUm3agN4cKD9Mxl7pIuROULwAUdWbUK
zHdy9aCYTIGId1IytlH3zba/xBB6xLz6gni0o9wsk0X9FSozvbC7w2/79hDx7YGRLzPpkq41hyFX4YJam3b6ly8z6ZKuNYchV+GCWpt2+pcxuQDwvIBSozEahw8xxHe+
T5akECED6hOtqvHfj1UQey8z6ZKuNYchV+GCWpt2+pcvM+mSrjWHIVfhglqbdvqXuAsVbJuXyWG2HI3RTClD0ijB45bpHUM4lW9Yc29yYoEePsXdHPrGiCaSEj9PpAI0
CKm3WDlS2yOAyORDRVL70wpJzuqvwwHUzVlz1AhLkcCJE7Q+PiUACXSIrCdNk1uMWzXU3PazDsKyEoFITyPF6m6A9aOVEKrrtfb9PUIf9qDy88crKpN65HKevWjV1A6B
CJGFNpzxBZQaBwzx706GkuSRSh/U1s4ejwV1imWTwknT8/06/U94y0/lzRK7DgOvcQqLIRRquG3rv23CdK3twEOFYCnYf6RbEuxfTq+igiYNFXWxON5rv6VTkvgZ9A5D
qVude4YVRSa1XUY8wT80QILEJGehoxOgc/jvDSGtKcb4OpUZGsPzPOdzn9RMRfVkf1XmWeKMuMWfg7yuQhFDZK1xJmjT9J0P3RaK59r4NOvKiCbRJr2HgYyrX3ljAm2I
KI6em2VK8rTntfzBS1o5AHoU0l8EMBvDotqDdivd7hvAQHC49OuaxebJZkWhm7drCW7CEm+W+X5QSwK8WKOd9uKbqT3Nzle/wIdeQdlwc1YIFrsHzk3H7lCvelokb6NP
N5q+XhL9gmVuQmR+a/eeXcoAprmd7vbLAVXg7FRctOLKiCbRJr2HgYyrX3ljAm2I3fDFC+1Zl/MG8QfQ7pbcYqEW36BOdur9I9q/kivSK7I9dt80r9szremAzZTOWVZ5
eCM9ixfVM5PEXOFC1nNB/1ScftTIYbW1Wfpg3KZqQyqGcbNE9qAOLEvcDkxFn6Qrrsqiuc7EFPdXt/CoU700zY+1qBcurW0bg0sSG8kogMCKBSWuAv5cpGLXPTOwMrBX
c4P2kONHgqskGsQRo59xxY+1qBcurW0bg0sSG8kogMApaEwYHu0PiB90f74HWx6rJLJAFV9g8hzr2FpnrvtKri6tPUHjei+LlOvuVQA6zjFEhaim2Wt9QpYPfnwyhHdy
eI5WiW7pKW04kkK2a/ONQIgo5nqny+DmDItt9IwXS9lTBg0XSc3hAXWjh0RAcJJgUFl/tkaIcrgdcBWeJDUk6noU0l8EMBvDotqDdivd7hvAQHC49OuaxebJZkWhm7dr
CW7CEm+W+X5QSwK8WKOd9hjURZKz9ALWatwhiDnQDDoIFrsHzk3H7lCvelokb6NPwC6SXHYPKxRIOeQ8ntsvssqIJtEmvYeBjKtfeWMCbYgc4KI6F8cpAJv6wJbrxhfS
taTW4dYFhcFEtLKogxAoejQr7KjWiXJ5k2G2lwIUfI9Kvzk1Gw8WKJQv9gSfjQ/k4yxyLl/l06g0ixpRTiLUbNmKN9dV4ZpyZWFPgbnl+uHbCNwKZQf6ab0E2f1jdinQ
LuJRNx4fyvAs4x7lKwLBAsqIJtEmvYeBjKtfeWMCbYi9wKHlaTnAw+7/GxBLn+3vzjvurGOaCzhIQUqtzs0xGliiM/UPb8MeEeONk3N2ya+UQyuB3ccr9idWeO5lJX9J
d8NwmncIGd+Jsa5PGV3rD8pkDWaFNJi4JKUghC3ej/mNuHybzCCVjbv0GSSWZ4QAj7WoFy6tbRuDSxIbySiAwBNtV9iR1jdMGTHrbJ1fwDTK2O3l/8k/5f0z1pUai6nn
j7WoFy6tbRuDSxIbySiAwABFMY50SBmF86+73PURyYE6J8K0PDDedHUMeYK9GKziN4be5KIleihjpumlIGVMmApwP5xLfuCkicxXIOhpxeMfsVQjw7rUAck03SNBRGSG
WKIz9Q9vwx4R442Tc3bJrwaXoQ2CHXS+62W9QdaKqjfeB6O5veC+wBClzvyIVV3NtaTW4dYFhcFEtLKogxAoejQr7KjWiXJ5k2G2lwIUfI9Kvzk1Gw8WKJQv9gSfjQ/k
4yxyLl/l06g0ixpRTiLUbOaoQJ/86NvmpoKGG50YO6V6kwZo/AEqx+IEuuWqYrkWWstj+K+E2UODW15yXBS5K72E9wv57flj8VPvQhXKMcxsayhHtedtOO1fUAYJI7rf
rt4WMfls2v0IR6labkuElw5rahz1W/QlnliBN8O3O/bMd3L1oJhMgYh3UjK2UffN0RZFXV7Bk2SAVih4LE271xXFdsdoz94eHkH/bkJZeUcKLRgqGtXfS4eDbSK/oTqK
yogm0Sa9h4GMq195YwJtiERYJ5VDynXSo4dOcX5VjJbcOQZYbFuwfQJmjgqLLIb9nH7t74/h4XSrPybIL+/vLZh0iXrC3MWeUoP9v9tb6m9paLCBfF+giq8EEYTqLGrn
bRJhH8GSN1DOAUhQGJLVcNC9tCyehhJfVmMkd0QKezCPtagXLq1tG4NLEhvJKIDA5cKJ1Q1MNScJN6BjQ/LAnWT5ifwr2JGmZX7TD+f7+1OPtagXLq1tG4NLEhvJKIDA
SmE0Q4DFQSR3jZb1WDWJfdc3aFpg9k6gdoo7/NWyu5KHdmrqBOulQZqhAKjxPWDC1JFvvIsaOz3ZZ84vhyVhNh54/X/5p6PBCQTzXYL4Yr7QvbQsnoYSX1ZjJHdECnsw
j7WoFy6tbRuDSxIbySiAwNW5/AVgI39wTkFnzwYdux5k+Yn8K9iRpmV+0w/n+/tTj7WoFy6tbRuDSxIbySiAwEphNEOAxUEkd42W9Vg1iX2EXu23fL+0MSSugXp9ONDQ
6AXH3jSKgw3oRVgK7uqIfF4fE3/e7A6i/M3Gw9VyEKXrnow0uUqrqaj2xO5jkCIanH7t74/h4XSrPybIL+/vLTEsT/u9CVVLBDC/RwPW5Q8GsJAHO954kg9+S+BfeAXG
bGsoR7XnbTjtX1AGCSO6367eFjH5bNr9CEepWm5LhJcOa2oc9Vv0JZ5YgTfDtzv2zHdy9aCYTIGId1IytlH3zUa+oP5zbsrKKChNoSzYfhwVxXbHaM/eHh5B/25CWXlH
35JhOV0WKrRzkv8nmbqqkisiTHFd2YcDiCnJeMGMknjTy3p3UH/oQN7PEZWhXJf7qJ84xwh43nQjZxhPBCL719v2yrZbIQCHY3y8nboRbUYezkZn5tvNf0LS7uuTmFIL
klPQVxw4Uhb05oAMZJT2IfetSo46JNIh2FMgyDkdWK6kUZZljHXeHHmH+uIEfS2Cyogm0Sa9h4GMq195YwJtiAzR8f7cttpbbNpFcpMUzQyIOg7YKkJtpz/W1itahaN4
MXelSorXtr3zdFgo3nwtaLrDPsa45hVxTBLWTpQaJJbiVxvsH5Kgg1xJDEWu/fYcoC+E5Dsy0uOcDbYup13Cnq/3uA6It9XuAR9HE2bPexOPtagXLq1tG4NLEhvJKIDA
0vHlt0v3+KOs5ro1ox4tdFy0o+izru9CbY2m/pBJDKGPtagXLq1tG4NLEhvJKIDAZ+j+FPXrK01AJDcfoGddh1NRPFOBwNEfn9/yT7OUJ9sMdNsVcyg6gmOmhpX83yij
VnSTJEdbmPmmJKDfEau2nxRMv2JgJtPzAC2nh9CquP8xd6VKite2vfN0WCjefC1oqj8oS2oVOAULntyWWrov2chuEZxgL4bQrkiC3+pQVycClBeZIAozHYwtYsdKrzfc
qJ84xwh43nQjZxhPBCL719v2yrZbIQCHY3y8nboRbUYezkZn5tvNf0LS7uuTmFILts1QXn0fBkiGe4ToMKIaEvetSo46JNIh2FMgyDkdWK7kazf+zIoLLD7TJobyxS5+
BrCQBzveeJIPfkvgX3gFxrvHqUY3pf/dTbXzfzGtbtkvSAWqomqOgzXJH2zeQ7HZWKIz9Q9vwx4R442Tc3bJrwPjzJB4N2HuBOfxOqogUpSxVNEZ+beOcqeICUhPubdX
s+rOB76DbYGn50lpAm8GwOXUhor+/mCFuGBpdPrm52day2P4r4TZQ4NbXnJcFLkraVnU0kpuEuTr47LzGTE5RcUP0NHEjciUsTvyUs2lxvmpW517hhVFJrVdRjzBPzRA
nsfqhqhJsQV03g7w6DPSal5gfdMKsIT5BEyiG1ArM6ez6s4HvoNtgafnSWkCbwbAUDXSu/xYDlyZVQb1mISnXI+1qBcurW0bg0sSG8kogMBOyE0/iBbQiCXOp6+5HNnc
lOfzE1JoEK8xPNPBGB5CaI+1qBcurW0bg0sSG8kogMCyg7K+KCsoLW4Os6mfpwbAWkAzOJMEc6udS4412BoFPZL7B3skzyV6V0aQohkOYQQFSxRDXTjMxYfvHxTkBbHm
tNzVmJtybeukxDeqjNx6D6lbnXuGFUUmtV1GPME/NEBujBhD4J7GJGvif0Q4GiG1S5ekHqOxbhFvOfXunYdzIDd2BlNW6XCsMWyal3NB4/8vSAWqomqOgzXJH2zeQ7HZ
WKIz9Q9vwx4R442Tc3bJrwPjzJB4N2HuBOfxOqogUpRwM3cJJ5uleO9Hs1HIRmvks+rOB76DbYGn50lpAm8GwEJnYCVrQExOyfuPPy+FWuo4QaZAOvsVW+kk/dOYU/lf
cisw6UJM5fl0Z+rctjRAmWljxRAE3Iq546RgmAjEm8Kcfu3vj+HhdKs/Jsgv7+8tFkgNHcjSGBBf2eJVjyJUfrd9WcZbFOTBoMp9sQAaO2WaIj3frYsws81ln2baUsNG
Ym7g4njev+mCxidod3fMkt+SYTldFiq0c5L/J5m6qpJmfZDuytXCrQ8Geix8wiQBZPLIxAB2VAzHIcjtUq3kj8BAcLj065rF5slmRaGbt2vdEkiKGd7RPow4mRiMHvkE
HCOYYRlgN6CvXa/3eYmpUZoiPd+tizCzzWWfZtpSw0aodFOrMt+Yfpllvs3KyVztj7WoFy6tbRuDSxIbySiAwM8u41DrZL9xrG/J7D5tmV+y8j6Rk/sw+8X36dPyXjMl
j7WoFy6tbRuDSxIbySiAwCEcKctpIqpOxoU6RmfkgoMuWwasyi8Wkhx16dXmKIfaeCM9ixfVM5PEXOFC1nNB/xB6dn9ZwbqV4u/VmOe7VJKWlU5a5exUx4+11ecLoP0N
qHRTqzLfmH6ZZb7Nyslc7Y+1qBcurW0bg0sSG8kogMDPLuNQ62S/caxvyew+bZlfvoDvLl646pJY+Xuy3tBWFI+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKD
LlsGrMovFpIcdenV5iiH2ngjPYsX1TOTxFzhQtZzQf+/Ko+jfoee0ah3LtdsY3CBlpVOWuXsVMePtdXnC6D9DemBfLQC961SLb1W2fqDg90vM+mSrjWHIVfhglqbdvqX
LzPpkq41hyFX4YJam3b6l/7T8x2atgyFiKhmqDAPS8n5Z6oHSra44zVCirkMoQoAfo3VrFHGi/HYFI/mU4GKWi8z6ZKuNYchV+GCWpt2+pcvM+mSrjWHIVfhglqbdvqX
LUAROClJs3ga2rba11LeM4+1qBcurW0bg0sSG8kogMAd3HEUrSOFhSA5/2fB7VLgUeUc23ei9C924gXgrw08wY+1qBcurW0bg0sSG8kogMA8VXvZ6b9S00xxEYIKU6L9
uh6Zrvvv9cGFgme40Isi4e2oyFHvINKiLaxya+ARnlqKqVAUTg+7LlCOjsUKdTjngptM+NmdpGSrXeZPXT5g9Zx+7e+P4eF0qz8myC/v7y1kfLxmQQJWSg+dML/NIika
BrCQBzveeJIPfkvgX3gFxuEA8wXfyAlun1kUeEgmKgtd7ScA8YNNWfGqjlbe9koGnsfqhqhJsQV03g7w6DPSaqCS61h+cPLBUKx4LciYmGiL7/tLHUPSEUkiHtDAVJd7
93epE81Kc+PbUpzuywIcm8qIJtEmvYeBjKtfeWMCbYhmQYTq0zIYtrp2gMnU7C2cMXelSorXtr3zdFgo3nwtaMxcWhjg+HjdG+ZntdJejM44QaZAOvsVW+kk/dOYU/lf
UAY3WrAd3GFeQxt2hWgFMYQoRJX83/ODOhG/syW1mhJd7ScA8YNNWfGqjlbe9koGgsQkZ6GjE6Bz+O8NIa0pxn7hlz8opiIeAdyeHlOPvneOMFDvk8QYIBnLjEBA8+5n
YqtMmuOKAZl/xk6DrOmNGb5xpVV2PRGZHsDnGntBhlNd7ScA8YNNWfGqjlbe9koGgsQkZ6GjE6Bz+O8NIa0pxgZntasLxWaxj/I4QDH7oBuOMFDvk8QYIBnLjEBA8+5n
YqtMmuOKAZl/xk6DrOmNGaXFdQ7sbMXzEM1KF6eJ7WPjr+j5usfLNOV6Urq1/jyAMXelSorXtr3zdFgo3nwtaOIC+/rCh2xf14HV1SOUgmNX4xHqhvwWKzvK8sCuCVrL
WGdzqgCwedHZ1Y0EFw4hwITIF/lyHhKABdw5GnQRfWsGsJAHO954kg9+S+BfeAXGotre+2aEnX1ZrgUDv1sTc0q/OTUbDxYolC/2BJ+ND+TjLHIuX+XTqDSLGlFOItRs
go+Okag2vOvUD6Wq/niELnqTBmj8ASrH4gS65apiuRb3ziVRMAZKIMt5IMJCgfzk2/bKtlshAIdjfLyduhFtRh7ORmfm281/QtLu65OYUgsvAQhwZhLt3fuJSNdY+QTK
961Kjjok0iHYUyDIOR1YrvKdMWZjelDU+RO6494kIhLK2O3l/8k/5f0z1pUai6nnj7WoFy6tbRuDSxIbySiAwDzI0n/T2uFjh1Hl5VTL3L+jIYR+az62q0U7MNYnJl0o
j7WoFy6tbRuDSxIbySiAwPMFzS0KwpEVQkOn0lQ/es9Ndw6jmnJy/QafnIfRVt7VHJLQy4ajfC+VyeN/EZs7SP6GN0PN5aU/54N/V5dV5Ia6t5HmSeW69xE+4x/Qrpm6
iCjmeqfL4OYMi230jBdL2SBeCOS+ySoB1QxAVxs86/+9hPcL+e35Y/FT70IVyjHM3P6wkB6vaSbliNcwnb9++Fzzsg5NyAtJpOhm36VgeNSYdIl6wtzFnlKD/b/bW+pv
lruBEzfrQnSzi1Q4FAd7EGJu4OJ43r/pgsYnaHd3zJKDwEKdYuYwF2IQPeupWEgpZn2Q7srVwq0PBnosfMIkAf3gy5DV0wTvCbGxJ/K9w4tYojP1D2/DHhHjjZNzdsmv
P+acVscvLdQOuyyhiU6nQB9g5nOkEOp/md3uPge15wegfZHaqrm2vGGlGMmbRAxvjjBQ75PEGCAZy4xAQPPuZ1zzsg5NyAtJpOhm36VgeNQWSA0dyNIYEF/Z4lWPIlR+
0x/6KSD/jbIDxax1Q3ArLPG9Kqkoxg4HFe+4g8ZlLHTODOmOcS2AgWIptZgKPFZkjjBQ75PEGCAZy4xAQPPuZ1zzsg5NyAtJpOhm36VgeNQWSA0dyNIYEF/Z4lWPIlR+
LVsKrzZdrQgJoGTtk8sz5PG9Kqkoxg4HFe+4g8ZlLHTxvSqpKMYOBxXvuIPGZSx0miI9362LMLPNZZ9m2lLDRvOKgXnvsOOIO0lzwWAbqItYojP1D2/DHhHjjZNzdsmv
jrqFRiOgjHW/b6TIYR6fhiVhuqsQK4vU3ouU8jHcqwu6YoHVpJD5cdqdMj91W7A1AY+CGuUsJL5ZJNMN0OmIEyNkuNPFdLIzLzrJMvhkCODHhCnkOJ79KQNeCYx0oGqX
gsQkZ6GjE6Bz+O8NIa0pxnUt6G9cqRAMZtFhidm2dM1/VeZZ4oy4xZ+DvK5CEUNkxKzsd0grMi7A9Nc1YwXHRTQr7KjWiXJ5k2G2lwIUfI9Kvzk1Gw8WKJQv9gSfjQ/k
4yxyLl/l06g0ixpRTiLUbCHWOAsKzKr1xR+BfCgpbyrbCNwKZQf6ab0E2f1jdinQR2NvtQW7nCs4O8nPs6/X5ApJzuqvwwHUzVlz1AhLkcCJE7Q+PiUACXSIrCdNk1uM
jzPvCBKnFTOEuri8xELUZ67KornOxBT3V7fwqFO9NM2PtagXLq1tG4NLEhvJKIDAzlokkZ3bSHowciWw+4nVPxx9PME6Evtu6lASEL2Tax73OF6t23e0aOJ7c1l/p4vA
jumoQ9gYpHED5tSDooyjpTkB3yd4Vs9gUPWbkqknKDXMRmUy5R0uLdNSCiZ+66Lo86kf4hivVKaWTa1DJyn1MAwCVRKohu2Y2GqAHtzT26H76jB0XKTasgRWOT9xOXA1
dJXRCxm9ylLO73Tm++LVrngjPYsX1TOTxFzhQtZzQf9pPxR9KcejEQg4Yvjxc3hVY3IeX0xIAct3C+O/J6aLbVrm0S115SOKPOBrIj1FjSOsyRsF6YkIo7eiJgI7SdeY
rt4WMfls2v0IR6labkuEl18b5dSx+Q2MiDeXGT9i0YftlDksGf13XNH9Yr3Z3mBe0/iGfRJ+AGP1gsC9nk3vXP7ZIx8RcvUasg8Spy1qojX76jB0XKTasgRWOT9xOXA1
/xKVZtreaQx/tCmlzC6KXR7ORmfm281/QtLu65OYUguLlexbvaQmzXOqbEhcq/IMnRu+6k9KS/9uQT10PQ6gcgVrGKZXso3JW8FK5CSc45776jB0XKTasgRWOT9xOXA1
/xKVZtreaQx/tCmlzC6KXR7ORmfm281/QtLu65OYUgseHLlk4WOPOnCTQMwkoe7mnRu+6k9KS/9uQT10PQ6gcp0bvupPSkv/bkE9dD0OoHKgL4TkOzLS45wNti6nXcKe
SNQ+ij3SacI8MlyLHNrritPz/Tr9T3jLT+XNErsOA6+1GwaxsOd8UYYLe3DW79MxIKkkM1KLIodm0PJ3s1iX867eFjH5bNr9CEepWm5LhJdvwhIQZSe4GJF/zkXNQngH
Mg9Iw0DpvkRgZAbSmZme0royPBdci1ZfXJOJ5bSwJ0W6wz7GuOYVcUwS1k6UGiSWT2igKwYDQF0NJqmOL9u8yJ0bvupPSkv/bkE9dD0OoHJUnsRlrmp888RxDgLj7QZr
WzXU3PazDsKyEoFITyPF6t0SSIoZ3tE+jDiZGIwe+QRSu+cxyKUW/p4bx+kf/hCF8b0qqSjGDgcV77iDxmUsdJoiPd+tizCzzWWfZtpSw0aodFOrMt+Yfpllvs3KyVzt
j7WoFy6tbRuDSxIbySiAwM8u41DrZL9xrG/J7D5tmV8BwFyg42GbvSF5pBJfbviOj7WoFy6tbRuDSxIbySiAwCEcKctpIqpOxoU6RmfkgoMuWwasyi8Wkhx16dXmKIfa
eCM9ixfVM5PEXOFC1nNB/1et/MbPqA+wgMzoA0icOJeWlU5a5exUx4+11ecLoP0NqHRTqzLfmH6ZZb7Nyslc7Y+1qBcurW0bg0sSG8kogMDPLuNQ62S/caxvyew+bZlf
rW5hGVHO7i+fws2huOr9vY+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKDLlsGrMovFpIcdenV5iiH2ngjPYsX1TOTxFzhQtZzQf9m3Y3Ex2qGGZG4PYWpyh6Z
lpVOWuXsVMePtdXnC6D9DemBfLQC961SLb1W2fqDg90vM+mSrjWHIVfhglqbdvqXLzPpkq41hyFX4YJam3b6l/7T8x2atgyFiKhmqDAPS8lbmVoOxXXSKv7WPNJxRlef
LzPpkq41hyFX4YJam3b6ly8z6ZKuNYchV+GCWpt2+pdg0ae8B15nkav494au1jS7CknO6q/DAdTNWXPUCEuRwIkTtD4+JQAJdIisJ02TW4xCOv8vOJ6X9xNLR6uqNSdy
rsqiuc7EFPdXt/CoU700zY+1qBcurW0bg0sSG8kogMDOWiSRndtIejByJbD7idU/A+PMkHg3Ye4E5/E6qiBSlNfgw/HdxD4BOk4Y5spE/LUMprgblUcJtWXvbwgcQhAR
aOuu8VOQ8929QLyrxdXRVwpJzuqvwwHUzVlz1AhLkcCJE7Q+PiUACXSIrCdNk1uMHRii5XJaDbOcRSDg8Sqd9wpJzuqvwwHUzVlz1AhLkcAePsXdHPrGiCaSEj9PpAI0
MXelSorXtr3zdFgo3nwtaB7ORmfm281/QtLu65OYUgujpxTm8sIk8hAbvqKE03daPb7Yz8zp9bCOmya/TO5VJgLuG4Q0JIXWlVHfZyQSUlOsr1Bhs61vPAmPfhJ7ap1Y
rsqiuc7EFPdXt/CoU700zY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwIsKSIigVCZaoiG2vlP6ewQYrPIwv+c8/jH7lzLpXrs3
lXt4s4cgo9zgkMS4YgNxAyO/oO2jYAIadg2b4t+LwWuPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
xahLLXWX+S1JnW8ZZ8FFoFcQrjKoIilvjhKDdDWGMmmPtagXLq1tG4NLEhvJKIDAzM4nXcdE6ECvYzuMWziVIWX8yJfa/hy6HODNqBa4JO4kyMduDmyBzm2hST25G11U
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMApaEwYHu0PiB90f74HWx6rBHQmzuIcp3WMGLAj7QG8ocoDpkk6SXGRLQ9sLUqBGnC7SWZ6sIEYQdCAsr8m53Mt
rsqiuc7EFPdXt/CoU700zY+1qBcurW0bg0sSG8kogMBUhlQ6qxQzijL1gMUihcH//9n53WRn+0AYh4dxS7MqYS2SQkTqRAPEcCG2fmDsNLWPtagXLq1tG4NLEhvJKIDA
FCgp9v6knUdJR0mjkoCy5V3tJwDxg01Z8aqOVt72SgZ4IRjxn+KU47EvPW/hkcktZsO7zH+wx0BkvHhBp3N7zGEwd9q/o8IJ+TG0S8k/hGbY3wjaFyYHqD8rNdP+3Ihj
9h/3dnFgaDhBCTFQ955m6rUFWRtPY+VRi9xy/dg0E0rxe/3CPqT1K2AcY0bkjANgzlokkZ3bSHowciWw+4nVP+tFsN+0jYFejjhcudnQYKC4JnfkZ0s9i+kCDYKUVx8Q
lDQS5T36lBxXxc5UMkr9OIlgLXrPGCyMjwkMshCrm56TewsVKdZXWRwPeNXPuD9m5QsBW5rmUWijN+QJvWS1gTvWEou3hju/2rdk9litmxRQebgaNhYZgcAH9lGP1F8r
5dSGiv7+YIW4YGl0+ubnZ6yoawn2+zX5AuepHsuLiAS4JnfkZ0s9i+kCDYKUVx8QzOBR5YRnrWFJuoQzsA3WgolgLXrPGCyMjwkMshCrm56TewsVKdZXWRwPeNXPuD9m
da6ztn9jYV46asZSyeaOIm26H/Nk2n0qxp7JF15iQT44C3VoPRgOEgJx6wxayTmq/ilmJ0vCD6QbjQS4Vo1FupCykMJBXQzcPobvYGqHm0wkrrC6etvJligNVZG3IKB0
AOQIFhlr3z4x84z0mgi5fyyuxQtlLGy9AydbHm+SB6sBj4Ia5Swkvlkk0w3Q6YgTOEGmQDr7FVvpJP3TmFP5X+ErJgYlMUMKU10Wvt+HFTYuncC6NqVW3xgdRCKWoQOB
Q/E5b0zRGqyMiB7cEtk5KrS4IKvmFrSZpI2sHO+R40e7yogS0VCTMEXfP3sdZDG8rOQmjJv4PJftTgvYtvgtj7SxM55/chSQKhqcaA4qP1z6s4g6X25FCM1OiMq9cJWd
2/bKtlshAIdjfLyduhFtRj9St9fpEL1Yq9FzO+MfiZXOv1sgMBa9Z4tzSh3fWyRpIN4z/ruvGyRyegvfb++QV60Xt71K6Gro+H2n7fYJS7L8CvFL9nXrqXZvAioIb0/7
KOyMzFEN3sdK/yti1qIvFpM5VV5JLUlaDj5yJOJSuQQZN8Q+y5nGQunpfb77fxjtlJr1aJ+p2yQkBHKmHxaUyLPqzge+g22Bp+dJaQJvBsCQsuoNBMFG2d3S+MfcyTVO
NCvsqNaJcnmTYbaXAhR8j44wUO+TxBggGcuMQEDz7mfxAaGhcIpBoW7FtOvY+1dvGX5ykc414Za3f6aqIzmbRQHE7xfIMKKDCpigK7+ZtPABxO8XyDCigwqYoCu/mbTw
VIJxgPtIZmBdaxo/Gxdjd5JaGHfeBF2T7ofFcCswPDAJxTvSUS2CGqdcT6nOHOTWu8qIEtFQkzBF3z97HWQxvKmOo2qdXUHSlXtTXp6dpoaN/1Pm1GdqYjRObP86lzsQ
Pu78FcypqKl3lTijVYVtG7vKiBLRUJMwRd8/ex1kMbzc/ICX3Z+x1RUvRC+RtQzVjf9T5tRnamI0Tmz/Opc7EJP3BDlr/nvSTeyT8s5WgoG7yogS0VCTMEXfP3sdZDG8
QxvdQoWsLxJu9tsNWFXml43/U+bUZ2piNE5s/zqXOxDm8xhF37QsxUSzMZuiSxARu8qIEtFQkzBF3z97HWQxvINvFkJMVDsRqDerrRYJaC2xuNuZfpH6yvXceByu0Nyh
8aWu9W9n7/PRNcJNqrbyS2kBf1Evh72MzG0jGcqym9lbNdTc9rMOwrISgUhPI8XqyjR9Hujryjgk9M9nZcmnoR11CJH8I5unnAf4ar76fO7jiiS7owNCuKhbmmRVE45P
V8BLo/8YJjPf1LZvaips+JVdbEEoNVIirzpiBIwH1ziR/7M0/YPm3Gdj6JPYm++bjf9T5tRnamI0Tmz/Opc7EIjaWvLLjlgrweez7PrJRbi0OA6YAXvQTo2U7B1BBRnm
yErGxGzU6h+jqPuQuTNkKxAKl/E68XL1kFProT6f4+Bkl3JiI7q1HhvuP73XQiylPRwDyOFLmd8B6yx27rw6LRX/RM3MPi6yuzjMwJURnBczLUc2tJ3NthZWZOLT0feu
1d6JlEeD2G6sNbXIQ5zFFQGPghrlLCS+WSTTDdDpiBO3r4LdpIkc4Vg5+v0nMt/jGWq850tqexZH+TsxOEJIT3EmFS3DCIQ6AdWTnDQVcgDVix1l0CxV2JZU4qIJVcRG
cfJKj17D8b+VEFIuO79Lm0ys4e5TKvVRx+CAm5tU/400K+yo1olyeZNhtpcCFHyPEoYIKzy/3KTGjITOBM4gCzSYzkrTR56TR20KP6ipILsq2xS1/K4CkswnmomrQq9n
NCvsqNaJcnmTYbaXAhR8j44wUO+TxBggGcuMQEDz7mfxAaGhcIpBoW7FtOvY+1dvYMblV7ETA71aFv7pNXKB9o9DxaY+qJ+pyPd/57+R2b2g96O5ZNtO+Zr0ePRhXDnp
S8fMFuamUYnF7jGGHi6okVs11Nz2sw7CshKBSE8jxeoJbsISb5b5flBLArxYo532WmKgU2pSHfPKAe4GgESNOkPQr18vJDD3nOZY7ZrCIOSOMFDvk8QYIBnLjEBA8+5n
YqtMmuOKAZl/xk6DrOmNGQF73dW0tNzgnG3tgr2p2tfe2DfolkiNM3wPtVD1H9WyT+g5CkQ/X9LiZcC5/9GwLrB+ZZRydMPWckrpFFKtSqFc87IOTcgLSaToZt+lYHjU
VTdN6x6a8j7oR0PclSiXv/PwWK8PPviL5Uz/X78dhMn8E+tNBjVDlHLtem6CpdNlIfptjvPa+jm0Pwxmj8LJIWNyHl9MSAHLdwvjvyemi22Of57197C0MhnxYZApP9v0
qVude4YVRSa1XUY8wT80QGINaUbJrS4DrO6eOCY0IzPZO2U3vR82WTT893XDAFrSXPOyDk3IC0mk6GbfpWB41IPFykBQkeLc5PvMnJ5Xb+L8bdpKxCZuqhDZYlHCdw57
961Kjjok0iHYUyDIOR1YrvKdMWZjelDU+RO6494kIhLHHJ7yoFWOX5fwKcdIhv4ujbh8m8wglY279BkklmeEAI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwDQ4oeGm0fnHCXTYbnF5sBl4Fa0tOp5zU+jyb7nINhA/NsxponKrA0eUvOSD6rLjxCjB45bpHUM4lW9Yc29yYoGPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAVNidUIcrJg98oXQz3EOw1fwI2kWcUTl8kNpg7PbByJq5ZG/yOfI37j5eX6Dbd1rG4ZE88BNAK01OxQxf8KG6x
rsqiuc7EFPdXt/CoU700zY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwAS+cQHqY3eFqv60vXHGV1WPtagXLq1tG4NLEhvJKIDA
MjFQIdAa/mBch1islV9uVaCJCM9mKoUjq4NumjWTnlMF8BUfn5g2NGIt41LSxlZXj7WoFy6tbRuDSxIbySiAwG5EHYsBkgPzrkYn+xFuyCMJJ4zO3pHkfusKaNavN4GN
j7WoFy6tbRuDSxIbySiAwB3iBscbxtpVTang4aPXCEiaUwXghaXt0dqac52xVDHhj7WoFy6tbRuDSxIbySiAwCEcKctpIqpOxoU6RmfkgoMJfEEAYMwBL0TBwfaj0d4C
DB8uSSmw7g7VoiSMRtWo2l3tJwDxg01Z8aqOVt72SgbTRr3fG1o+Svm/uZXL7SPA7Nk8YZ9j2UKogLIFbTsDl8cp8UR1ywOtnbZ2c0OxBvcAjPNiQ97jOo7wV4PS92HT
iyQcxxKZ6G4H5Pqg6MnfHOZnwW/4X4fux/9uvDqubOVhi9FYkvwtqdjEP55SEUxSgU+F5smR0PDar73OhYjlbo+1qBcurW0bg0sSG8kogMAd4gbHG8baVU2p4OGj1whI
ZKswxd1bzN6xrvvGzJvdl4+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKDCXxBAGDMAS9EwcH2o9HeAgwfLkkpsO4O1aIkjEbVqNpd7ScA8YNNWfGqjlbe9koG
00a93xtaPkr5v7mVy+0jwHyKvi42cj9aUZ5PzoTm6LPHKfFEdcsDrZ22dnNDsQb3AIzzYkPe4zqO8FeD0vdh04skHMcSmehuB+T6oOjJ3xzmZ8Fv+F+H7sf/brw6rmzl
YYvRWJL8LanYxD+eUhFMUoFPhebJkdDw2q+9zoWI5W6PtagXLq1tG4NLEhvJKIDAHeIGxxvG2lVNqeDho9cISIPEH7oyrmdi6nmR8WcwEWiPtagXLq1tG4NLEhvJKIDA
IRwpy2kiqk7GhTpGZ+SCgwl8QQBgzAEvRMHB9qPR3gIMHy5JKbDuDtWiJIxG1ajaXe0nAPGDTVnxqo5W3vZKBtNGvd8bWj5K+b+5lcvtI8Ds2Txhn2PZQqiAsgVtOwOX
xynxRHXLA62dtnZzQ7EG9wCM82JD3uM6jvBXg9L3YdOLJBzHEpnobgfk+qDoyd8cx6e5K2f+0/KOWAbuiisQgmGL0ViS/C2p2MQ/nlIRTFKBT4XmyZHQ8Nqvvc6FiOVu
j7WoFy6tbRuDSxIbySiAwB3iBscbxtpVTang4aPXCEjG3tWNsZ757ggdKUSkx9Tkj7WoFy6tbRuDSxIbySiAwCEcKctpIqpOxoU6RmfkgoMuWwasyi8Wkhx16dXmKIfa
weLX5Sb/SBc/N4s1QBMXrE55cZPYR+JBWgefKC/4O0SNuHybzCCVjbv0GSSWZ4QAj7WoFy6tbRuDSxIbySiAwINn3C2V6q9OTumJqlGyb4aNuHybzCCVjbv0GSSWZ4QA
j7WoFy6tbRuDSxIbySiAwJ5Xsv5RaiqkXLmn3hFKLaKybMfgLQSh2U9GRWe9/5QAYfJffD1YNMST4aW+FKT9woskHMcSmehuB+T6oOjJ3xzukiGgoDzdjjSs2n3pdbL6
YYvRWJL8LanYxD+eUhFMUrkYgGA50ec4iWZjwzhEgIRh2gc7eGvIMt9Vsb7oTM9BcYCOiAOxQ6y7GnoG12rV8FL7NE2xxFQIceI60pt4YXLKZA1mhTSYuCSlIIQt3o/5
jbh8m8wglY279BkklmeEAI+1qBcurW0bg0sSG8kogMAhbhZOZzMrsKy/RCj+Fdltjbh8m8wglY279BkklmeEAI+1qBcurW0bg0sSG8kogMCeV7L+UWoqpFy5p94RSi2i
F5T5fP+45evJnB/X2nkKZHesMdHzVDlGVaABH3rgs4kh7JQtj6ONZV2j4lTwOksXj7WoFy6tbRuDSxIbySiAwEFEapOafIXnyqUwCLo+PJi9u8XwNrdI5932YnJDpUam
9hNoH0iJDZnuecE30s8yP4+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKDCXxBAGDMAS9EwcH2o9HeAgwfLkkpsO4O1aIkjEbVqNpd7ScA8YNNWfGqjlbe9koG
00a93xtaPkr5v7mVy+0jwHyKvi42cj9aUZ5PzoTm6LPHKfFEdcsDrZ22dnNDsQb3AIzzYkPe4zqO8FeD0vdh04skHMcSmehuB+T6oOjJ3xz6aDE38IMmUkj+D2oD7JBq
YYvRWJL8LanYxD+eUhFMUp946hB6BbxjIXw2WI5PjGWDsvK+/Jt0twIy5NnLF+VGKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwBU2J1QhysmD3yhdDPcQ7DU2unVc7bwUz8QQEi6CGnRYq07JqQqbS611cpFK5R02Rj/K4GDq7kQ/vViRN6CZ+0qPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAMMkpQWA3gtEODlAoUS6V8o24fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDA
Wf5s0PuxtgTUL8+pRYJYziPvL5eNdRgnZzDO89YzdKO3oQqQQsWBC+z+zmo/sctHj7WoFy6tbRuDSxIbySiAwIkTtD4+JQAJdIisJ02TW4xbNdTc9rMOwrISgUhPI8Xq
69IRjaJAPq+EPYzwMG1wMKM/q/uOQI55PPS278oTGzKyaSZqX63L0ZQRSlf4E6iFj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAOJeNJZZNPvfoOAGtB8cJW
21urzb87Rqacwd1UZGRuNVcQrjKoIilvjhKDdDWGMmmPtagXLq1tG4NLEhvJKIDAzM4nXcdE6ECvYzuMWziVIeeCTjsKmV+/vwuRRUrb7OrLMhpYq44Yk7QVSYzxGPhA
nH7t74/h4XSrPybIL+/vLevSEY2iQD6vhD2M8DBtcDBy5w+6/PeV9lrFxsHsfBlyjn+e9fewtDIZ8WGQKT/b9KlbnXuGFUUmtV1GPME/NECAw0xbb1YIeDQBVRWh4td1
OCOphLsjoh2zywQoi5XE42Ju4OJ43r/pgsYnaHd3zJJPBn1jsatS59Q2NIjGnl3MKMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwPf0yNZJeURuGK2os6GGN7D3Xahj+AvJZpN16PBcUpaGjbh8m8wglY279BkklmeEAI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwAaDiVsCDvQgwfmHf0imfy7dxvKh9ZMhw/36feIv7oOkzMP4PUjGHbsd2A8mwsaKrohYAB9m8ojGsmFrWLKm8idzg/aQ40eCqyQaxBGjn3HF
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAYzo7S+/XGUYuj9JQn3nuYy9TC+PVR7Ebe+C8+bq23EGPtagXLq1tG4NLEhvJKIDA
Hj7F3Rz6xogmkhI/T6QCNP7K1+bpJmsDvZZ0Syxjnsd63xvi6GlEUJknxEfSAgvtCknO6q/DAdTNWXPUCEuRwI+1qBcurW0bg0sSG8kogMBKYTRDgMVBJHeNlvVYNYl9
0F/5g2oWbB868H7fU5n9vovH9BXI9w47FB3KaqIVq/sgSYyvVtufLF5ns0ScUSSMc4P2kONHgqskGsQRo59xxY+1qBcurW0bg0sSG8kogMC74w4wEBAepOCiQ0nq3dzK
cEARDUwEm7/5ltO3u7bFMckEQGAgtrNvMUgEDrrXfR2PtagXLq1tG4NLEhvJKIDAHj7F3Rz6xogmkhI/T6QCNDF3pUqK17a983RYKN58LWirRPhm3NZJzoTYvk3gDjhJ
mb8ouV4VrvicSGSvYjqG92O1HlOqyNaNYPeOJQ+5e3DF5DbIE/zgLmYt6wl6VNSygM8TSanF4ePTFFuTSd/iw2N24MOKqLPOd/OoIYsvt/qdG77qT0pL/25BPXQ9DqBy
JlbBrmIIO0SKWQQtLg6EkLFI2PpQuPh+cOMSlGYdHJo2nSUXsvnVkBSju2V+3ojpK3DruWJ8Dj6GeBWZH6MCiFPlwrykyYY4NpYfbgWibdX2NCqPGaL52Cxoarg7W5Py
y1z6FPksj/zp0GY6Vu//4oSm2O6KJxGWPfGe8Sx2+jiHBohUadBw8UXgfGqKtwijyogm0Sa9h4GMq195YwJtiB4vNDHFbjw2lpA/nYqkjGe6ZK7+yzlQeiQAc6yh+zEg
mukAWE2jZv4tEmLBkBSFRJYj6leqeInqYSNsaqoK1yr35Qqp600qBxqEyT4mgDqQDUKyAKr+JHgN+lvIdEX5UWc3dRclwJRsEyFcKtPSntha91jsvZr1DNI/1jRBgCVB
9W/XftCUaKQIplwKlYJToKTrHBeO0hlALBiFUSlQ3AKTZR1rQkLnXHTaTy4J1fJxK2isaj1BtXkcGgF6CEzrrv0vfoZLdHZHkUTjL3TwKg3lWYBedD6hFeKSBRyP7J0q
OzJJEXp+33mcMGDK6UekuTF3pUqK17a983RYKN58LWjtlSRrVKKC5O+vPdu5vF9HUrXZjqacw9D/OeJZYOAJUrwpvm97BH2mdJUBOY0d/150vv4ch/Gi5439gNetQ0g7
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAL71iCCWp2Yai5SbdqA3hwr/4RziVJYLj79C+iQ1toEjangJSUGxXx/UwjQU6GR4g
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAGeaCSKLJtqBzjaG27/0ZBE+w5QjoOrBFzwjKa0tqg8IKOBmPFO8XIrYVOs5kk6Up
SdKBsk3i6sNPuyXhUkIx0I24fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMBlwzIuuC4GmF0cXD1Mx338
3e9WGUAvHXVRNEr0qrBB6I+1qBcurW0bg0sSG8kogMCJE7Q+PiUACXSIrCdNk1uM8WHpNE8KWS6EvFj2bY6o2lKSx0bueFI4/TLTOfFX/JyuyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwHhunupN7vLvEaRZOLQP1Zwp/ebEKxJ60OVFLJpTERcvahuGHWABwh2Hq9auA/2eRSBJjK9W258sXmezRJxRJIxzg/aQ40eCqyQaxBGjn3HF
j7WoFy6tbRuDSxIbySiAwLvjDjAQEB6k4KJDSerd3MpwQBENTASbv/mW07e7tsUxyQRAYCC2s28xSAQOutd9HY+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0
MXelSorXtr3zdFgo3nwtaPxH3+n3vWaUPO49NEjDfJ3mS/i9C7BoGvy/PaBQVlWYWKIz9Q9vwx4R442Tc3bJr+pmjhTtWAYHyGn/IMsvvFcSybHBd0BeUvU3NYE+h1hc
MR1EmMuP/5Zl7qxkS5cvtOufQStaHEUs/3xZ5ASoqMeaIj3frYsws81ln2baUsNGYm7g4njev+mCxidod3fMkgqCkuBj0f9GZthy7Rl8ZZH1JzTPktUdeeBwzGSXrQgJ
DpGrrv35E9NCANKWf7hjDbPqzge+g22Bp+dJaQJvBsBQvt1dgBka/13BhGVOoZICCknO6q/DAdTNWXPUCEuRwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwBOgJeHxYFzLopWEdfTcvCGO5QUVTZjZFYew+TIAwGUVRm0DeqRi7Fc3T7azVeVRZ4+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMA/64XqD7O6lLtgbDnzfQxYcuho3uW3qzsGw5yNdIECzQwtgm3/lcpeD1Ec/5jOOQLZ4YrvKefB4NEIbowBJ4Dq
KMHjlukdQziVb1hzb3JigY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwCAdsX5+3glnHjcjW+zf/T7nL6UdBtRtat0THdyTWKMq
j7WoFy6tbRuDSxIbySiAwCEcKctpIqpOxoU6RmfkgoNuAixn85A4OSjqFBWyMOl35AOKcOfuOE/35xJ/ri/67o+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
nley/lFqKqRcuafeEUotouODkmCRQDPaDEpUM5dH3jSMneEnvBcEBU3ntQD6+O+Gu0lmerCBGEHQgLK/JudzLa7KornOxBT3V7fwqFO9NM2PtagXLq1tG4NLEhvJKIDA
VIZUOqsUM4oy9YDFIoXB///Z+d1kZ/tAGIeHcUuzKmEtkkJE6kQDxHAhtn5g7DS1j7WoFy6tbRuDSxIbySiAwBQoKfb+pJ1HSUdJo5KAsuVd7ScA8YNNWfGqjlbe9koG
IQhCRZwh/aA4opgC9EwsjAqNHa0LBKyQ9ZIMuJZzlDOCgLZVCmpARKwpy4CBIxGxiWAtes8YLIyPCQyyEKubnnJpHf0Kk4RaA1Aobaoxq1GYTyi1OS27lz7KS+CBexzX
YdoHO3hryDLfVbG+6EzPQSXJr67GnbpL54nvPbARsXM8Qf+IoWy4CKZWveGvm45UAcTvF8gwooMKmKArv5m08Ir9Z8Dluws3C+RAa17xDhPAQHC49OuaxebJZkWhm7dr
Lv48jDwLuXWtHY/ThAbd9nlerNRo96dhXznteoL3PaGgL4TkOzLS45wNti6nXcKeX7OC1f3ENmYJfDc8UjLRY4+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMD4V5ByGvSX83epI/kjojqmNVOxDEsYVvB/WOwCakgqHuw8QLX6DdJ4a9fIlCwNbs6PtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMBX/H3xpUBTMW0mYSoD9oQmOQOzAmz475ifNJaVYrVca1OOxesHc3O65Wm0Q/fTEkmAMmMQ0uSjcveIZs1Fjk64
TOyQLELykG1Z4QoK2E0FxdPBU0kfhE7N9/sfmh+uc1WSqy/0JwXnrgxh9PHca+yrOn3cVy6Wm6Be14gwZxliyLYlln4o0o6SpqAAE0s3hBXjD/te8gyoZSXpe7D4oEoc
MnsLtn5PK3EdIvoNZ0jxPy/gEz9vRqfc0ORnapHijUCGk8qLdeyoCJIlQZNkpA3us8J2fmX4jlMjDdAa8mN+Fo+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwCQ3iDsa26VCbi7qBViwuHcoweOW6R1DOJVvWHNvcmKBHj7F3Rz6xogmkhI/T6QCNGa/vj6NkxvQMwCbp9I+zQwF8BUfn5g2NGIt41LSxlZX
j7WoFy6tbRuDSxIbySiAwOoYcxaJt+VUCal+VeCKf6p3mlPGzc8Qf7RrKwKsE7cmj7WoFy6tbRuDSxIbySiAwI8qeMp9yQj4gifY2gYG3nIfn0/yKyjQ3YMiXZVaI8JK
Gcl1gDEO1xjax2hiiG83Lo+1qBcurW0bg0sSG8kogMAwR/1lic4GsBlki3Qv5fGOKu1FlsKYb3L/jy+XzdGkP4+1qBcurW0bg0sSG8kogMDPLuNQ62S/caxvyew+bZlf
kARby61TZfxSoXJxn9rP84+1qBcurW0bg0sSG8kogMDMziddx0ToQK9jO4xbOJUhcRKygVIp/4M/GIBbsFdDM06AWxn+8VfvRr9gP58LTm0sccJIh7/IF4MO3CzltN6J
8gJ49+TSnK3f/G9NcJvTcggJ44gZnViodYvoqebYWEKpW517hhVFJrVdRjzBPzRAks+tgt0z37/ucubtH7x/A46FBYfQd31o6QKKsLwIv5Lb9sq2WyEAh2N8vJ26EW1G
f1blLSfr1oVDtGioS51OdVGxZ+5RbcEOAF/bxrX2fD7n6KFdPYgIPlYUqXFW45IyYm7g4njev+mCxidod3fMkvOKgXnvsOOIO0lzwWAbqItd7ScA8YNNWfGqjlbe9koG
+UkUP0rIpkfSwq+yX8yRsB26LQodE499Pj+GJaT5ebZJ6VJOqRs+16UgJsZsetG+/wCw8Z9KwwNpYlpQeXe/v50bvupPSkv/bkE9dD0OoHJLx8wW5qZRicXuMYYeLqiR
T43SoaEPYNNSHPwwJ4jlvPBN8ZUuEMNUKXbi+DsVVSeIRmsED1sU3EWdzpvCXeQThnGzRPagDixL3A5MRZ+kK67KornOxBT3V7fwqFO9NM2PtagXLq1tG4NLEhvJKIDA
hbKo6VnO/7vRNfddIfip+q7KornOxBT3V7fwqFO9NM2PtagXLq1tG4NLEhvJKIDAzlokkZ3bSHowciWw+4nVPw8iYnEIgkZfeU5e9RMv6wSi/niHH+i63aU9MNiU2BX3
yG55VjyZKFwgWiumreBq7gzEIdoWQ6rkKpIlu1o5b9OYREn4q8YJxeRQ/qeeSulMaa6Hlxh9queHjDDvMvv1KX9W5S0n69aFQ7RoqEudTnXwPJaKGU6LNSVR+YhPovz3
iv1nwOW7CzcL5EBrXvEOE8BAcLj065rF5slmRaGbt2vkZc/3S96VbJQflld2YiGM4NucbS4Z3RLnk+usiIazeJ0bvupPSkv/bkE9dD0OoHIh7JQtj6ONZV2j4lTwOksX
j7WoFy6tbRuDSxIbySiAwEiLwFB/2qE8KNs5e+sT6HXqjWcxwyWbZnTwZ9fkUAPcj7WoFy6tbRuDSxIbySiAwLKDsr4oKygtbg6zqZ+nBsCJtE1CFZPyVQbU8Gv+1nN1
WtaxtPjsG7qiYbCqX0IbzPRrd9AjlpGDPE/w4OSCgTOw2DmMEqVuEhwyHzykNCMvlOlDh/1CdcsupVSce59jYNPz/Tr9T3jLT+XNErsOA69Zn+iFzv1LIZe8gsY2G1QW
WKIz9Q9vwx4R442Tc3bJrzPJwyE0zJ3Klk76qky2pTc/M4gAOXGRtaXqwOQIWAX4Nuav0DwxPG/KVa/UGzCNSbPqzge+g22Bp+dJaQJvBsCQ9V0PxO/jpKQxaFaXBMOK
8qZsxc2OgWpl/rVjREz6rdvnlwdVxmnjfKd0juPCaqyWP/+loT2YQKUUkuY3l9w/V7F7jVeVyRy2VkC9oWmWGlFwGKZaC/G1mlEekwCNiXlbNdTc9rMOwrISgUhPI8Xq
5GXP90velWyUH5ZXdmIhjJ3I9P4WTbvHfhM8FSggSY5Z+S5lbr98WCWExjTHNYdM4LzDSEvvbmCSudcuTPiwxP8AsPGfSsMDaWJaUHl3v78FaximV7KNyVvBSuQknOOe
wEBwuPTrmsXmyWZFoZu3a5ePJ9P5AkOam38wAj7RGRA4Cu8hD3baCUQK+3DJUjAUdJALm99oJlbWIUAK7CpzmJVdbEEoNVIirzpiBIwH1zhUnsRlrmp888RxDgLj7QZr
nH7t74/h4XSrPybIL+/vLSbjB47PbKnvX+3Xc5b/m8vpxBy1k0mjV3+4jRcYOOjW8p0xZmN6UNT5E7rj3iQiEsrY7eX/yT/l/TPWlRqLqeePtagXLq1tG4NLEhvJKIDA
Lbu3In7BeqLug8wUMipJjMrY7eX/yT/l/TPWlRqLqeePtagXLq1tG4NLEhvJKIDAAEUxjnRIGYXzr7vc9RHJgUpDTH2IA/D/UKR20rM2cM8fMU6XuUx5D+bjdHsRLn8M
OcOenTOK7EoDxC9fgvX4ezCawo7vgjgiCG02XO0zo6WPMb+MXOr4+fUdlu5UTtedcMjAt+NCBFMo4IqrgoVp2Z+X03wLglDJgIWNLQ+2VGSaIj3frYsws81ln2baUsNG
84qBee+w44g7SXPBYBuoi1iiM/UPb8MeEeONk3N2ya8jzaqdcUosgeUF09BWmhjUWKgxhNvj+ZNE+yaH8TyeACNrILY8hRbR8QDvlw3ypy9zg/aQ40eCqyQaxBGjn3HF
j7WoFy6tbRuDSxIbySiAwLuOMOlv70OSTZzKy0zApSpzg/aQ40eCqyQaxBGjn3HFj7WoFy6tbRuDSxIbySiAwCloTBge7Q+IH3R/vgdbHqvWwn45bHI7PoTwqLjQbxHR
viPBUfMABYZu2PJ9sFxgbDu23OaGruaHOX+YM8Sr1SfAQHC49OuaxebJZkWhm7dr5GXP90velWyUH5ZXdmIhjDLeKbljYbiphDZv2iyoF4edG77qT0pL/25BPXQ9DqBy
S8fMFuamUYnF7jGGHi6okU+N0qGhD2DTUhz8MCeI5bzwTfGVLhDDVCl24vg7FVUnoOLMlZyJn4W7dJ8OCsHi1IZxs0T2oA4sS9wOTEWfpCuuyqK5zsQU91e38KhTvTTN
j7WoFy6tbRuDSxIbySiAwAvIWukFlHt3+GtxoEhNub6uyqK5zsQU91e38KhTvTTNj7WoFy6tbRuDSxIbySiAwM5aJJGd20h6MHIlsPuJ1T/rmWMMil8a2XpEav4SWg0U
5NhzgySgqPd0rfWIffBLxcIvujQ3J2UHZ3sbpXqQrGgdBa80UpmsoOdd1lFNIqKs9Hv8v7VLcdMMPybouyQQFViiM/UPb8MeEeONk3N2ya8jzaqdcUosgeUF09BWmhjU
FY76DqgDwIR2k+9HR/HOj1oyxVfOdk5l+JXgqPeBxVyJYC16zxgsjI8JDLIQq5ue3veY+tLnIpqyWQwf38kvGBktOP/BVAM6p3ToB9YE7vCz6s4HvoNtgafnSWkCbwbA
UDXSu/xYDlyZVQb1mISnXI+1qBcurW0bg0sSG8kogMBFPS15PUqdWcFUrTh17GfFfpd8ist2RnMzzAJK74kvmi1bQ2BjJVjP8OQtNkHGTgiPtagXLq1tG4NLEhvJKIDA
L71iCCWp2Yai5SbdqA3hwqZbHdPt9hVzl9aP1h3lVIXyRU3wDUQlxyPj5ui/00OUXm44RJpr38JUdfIBPV+AOYjBCUIsIncJ0vpn7sLc3GOcfu3vj+HhdKs/Jsgv7+8t
JuMHjs9sqe9f7ddzlv+by+nEHLWTSaNXf7iNFxg46NakUZZljHXeHHmH+uIEfS2CjzG/jFzq+Pn1HZbuVE7XnXDIwLfjQgRTKOCKq4KFadmfl9N8C4JQyYCFjS0PtlRk
miI9362LMLPNZZ9m2lLDRjJuloTYVUmyWqKOD8i52hITLUfXC4yzvL86Dx9Z/93Uj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwA8yLaG9QZQ/ZK4Dv2bSjXtIGJU3FnAPmeonljiwChSTueByvdfN80B5F7EN0WeUCft0I5BeEGSEzbZ1oqbCtBKPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0QYJTd9igZVCwpndHvbhUGa7KornOxBT3V7fwqFO9NM2PtagXLq1tG4NLEhvJKIDA
VIZUOqsUM4oy9YDFIoXB/9GmRw4T70F4G+bXrz39bLAhlbkRQiLfck8HwdnUENWKj7WoFy6tbRuDSxIbySiAwBQoKfb+pJ1HSUdJo5KAsuVd7ScA8YNNWfGqjlbe9koG
KmLopWVHLXnBw3OGwId2fflCK2Dvux/4vZ24L0hx5123vTaBQMsJ7Uy0Cp8hvgvbj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMABFg5NyA1mlyMaKOYJCivA
KkaN+OEwxvPh2e5XbQ355424fJvMIJWNu/QZJJZnhACPtagXLq1tG4NLEhvJKIDAPFV72em/UtNMcRGCClOi/Ygo5nqny+DmDItt9IwXS9ml4j0NwvY/qEnJFRXZUK9O
JK6wunrbyZYoDVWRtyCgdHBoMkHTmwp/ug0j6avE37/lARFAOYsS+Gabp8xeE9ucwza0T+uKhY0BgOcgDzHpiUimEVJJczlFF5rrFqjO6m1PYcmIwHODUJie6wqz17kF
SyDJszfznQHE1H+eUjvs7SoY1joCIvMWP0xKFT8hTCCuyCcH3NKNi54OjWYgXTg5s6GpcMkEY4PKPMTSMXlMskXp7SeKVkqHSOMZ7KL6KaV4jEl+dz8MttzsfJPq1VaB
yogm0Sa9h4GMq195YwJtiGhH3yrAxZjo40083iog2Wxi72hO362rM3Ekd4COxVuhr+faAdOJZIRkP3ghpqvZqPh3Beh+ljmJzxNosek49HLeeflpwfYJqB9t2+SDbbZO
s0ZwWSR7tmK+7DD5yIm/CHe0qlpH16/JjNhQoOrDawn245dr/RhXxv5XW8/Og/7JPXbfNK/bM63pgM2UzllWeVgUA5ZkQsfWunll+6/shkrnJAFRTAU17kfLPUE13fRy
VJ7EZa5qfPPEcQ4C4+0Ga5x+7e+P4eF0qz8myC/v7y1bfV73/pMt968X1Uw8fRRvPavesGxz3bEYNMkT7SuGRfKdMWZjelDU+RO6494kIhKodFOrMt+Yfpllvs3KyVzt
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAiRO0Pj4lAAl0iKwnTZNbjGu7x3Qv1Go1PUinzX1CzoD6Rlf35k0Ox45mQd0X+3TD
TVw9Yy0dUDxhaP0IXY9UvY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwBQoKfb+pJ1HSUdJo5KAsuX+eveHbn2p2Y2bcXssPquS
Jpu67XpGdbRQemxKameREzCyQvn2T0voOYKV60kGy7c3Kt7+vSynYOXH+Uu557GCtE5q27p4jv3wi2X9Us0J4Lzfsr/LT3dHeXbzACheC6uG0mdWYHbHeRkCxkLItbEh
f5lgpQAhD+P/fFW86ULoZ3/nupP0Q9FecdSjz8crlGRnyosbpdSxhHxRw8QRcDAIyogm0Sa9h4GMq195YwJtiJ21V6q5UBlDxG/RkYAFJpzMvSrpg15PAiZ8UdzbmxaN
8SiKUUs/dfon8XwXlCk7LQyE7GUECOQMXUerCd0NJV5xkP3QUhx5AooQf3JfpcT4ueEr5ncQOEBO0RZGYiMkw4/BS0CzJVkT73VlWfhxyjGOMFDvk8QYIBnLjEBA8+5n
J20TSj/4gQAb6YYmWdIWKlUxxednYwgBs3Q7KY/tE0+VvpNSmef0lYHyPebyZOaRQ8RO4U30EIDayscVzIaKLo4wUO+TxBggGcuMQEDz7mcnbRNKP/iBABvphiZZ0hYq
aQEzspv5UfPbgz43BDjNWbt0LwFGH6YUOeLkrjvow8c2hTOA2HRSjkN3PcYPb2dLyogm0Sa9h4GMq195YwJtiHcbERSzpX9dFNTmfyvupHOc1FmcMtgJfQpOMHS808sm
vvriPb23QQQg9HYzPAtZR4WJ0M7q4e0mQI9LTLRRIA/KiCbRJr2HgYyrX3ljAm2IdxsRFLOlf10U1OZ/K+6kcyTl0LMdmu/FXXKPfM8pW6CLF+uQ6zM2fOsfO49HfQ4z
k6orUhQ/F6Qc9FUKuGwhDcqIJtEmvYeBjKtfeWMCbYicNTAIxNxV8BpoP51RVXG4nQuT66BfQBy2G+JyNO4FlxiJ82XOKt6iNmtyF8qKrymrpAuOXRpkdIsvatOqykCJ
yogm0Sa9h4GMq195YwJtiEuu2frbXRY+1WXKvIEH1JPKiCbRJr2HgYyrX3ljAm2IBqBwDcEy5WCaUWdM4KQfFtcJWWUb/7xtGqeU3GOwKa3hHBG9UkNDVkKhPlVJ+Q5P
q8jYn8t1QS6KWD5N533MtzErQaab6iRt33Ev+5hlJYoXzle0e+l24QrC9GtFg7f2g8wto/vu5ltYfmLdC1MVU8By4efZTHffq42g9ZnjF8pdTGsZrjhM944etSsIRk/D
3UHfZitakH7e536fLub9CbMAO7y5j99aCUNSDQZRLAlYTicCCMm5myIPHm4xZXjwY1bf/xnkUC82GyomZkpN6UhcFl8BO7vz3Br1UajwEzVof9zlsuz1ZOOpoQLnapfp
g8nm3e3/Vq1BWRI+x0XVdoYA/Bq0DBNaeH7SU+aU/aFU2LIMXGfHe2cSbe9pW1Z0niZOj2bxCVKef0bwtI26ziCTtHHAHZUw3eEE4oZOfWWqsAvnj3OITMGByP/j7iIZ
A+pt3Lg0FieYNfrST0+8+8b5b3xgl2x6putXHoOrkIPKArBRpT6RZiUBRgeT4tk1peVftOdY6ZPUflWnyeHena82ajNi1pn9qROBeOH2HyJQcGit7VzDiua8BHy9Ic7W
CT9/iS+mFUhpHugnw/XxWJGBZ7uAuW5E+IpTC2P+mHjLyVfc44fC1VDUwqTANhHvoEl3IYtE4MaA7CrhqTLIz2s6AbnZPBUqCp+w3MBx8YOLjSzInPZcuwbFPD3RGRPS
cu7lSCf6kOEYJJmqjiv3p9bHwpY/jWBoBTf6TwhuxLePtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMAePsXdHPrGiCaSEj9PpAI0
MQPKegienInrQ/N1cWBrtCrisIfrBar7U8V1YYHt5qgKSc7qr8MB1M1Zc9QIS5HAj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
q0Zm4wZLCvH62A1iGN00W/tYQxGhVZdUqT21oFvStJmkYkb9hGj83Zz1ixh5rMkxFXKt3DsYIJOqhsLjS02UaE6ICDeIgVNsk8IZSYoe4gAc26Llo41jIH/a3Bxg9uHl
QYMlkRPcO+wkoKwThRa2VgWBszCCjqJoY6DmDAxH7uK3v+uYpbsIyGXrshs1mrS/cEUFRW0n2MZy5LramiCYJ+h9IthylWEmrHW63ViTK0zvBT2P/kAaDAQ4utR8tGFo
rwNOhx17bVCyOhckwGfLcNPr+A83KXvN7QpJxBSADXoBhqsQT92pwRQfnPqziOoaj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwOwYDgwLjgwfDLdUCmRqIZIshg0fhQrcDafuvzHIq1mXlQstqPRm69ySx+OqV8elyQpJzuqvwwHUzVlz1AhLkcCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMDgnO8cX1xGleIeJJIAQp1tJIs5czDUlGl2tde5POsoRk4zCL/ggVDncwk4pbLUfZ8Q5vymcv/QHYhFoXMLwt0G
c4P2kONHgqskGsQRo59xxY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwGM6O0vv1xlGLo/SUJ957mMvUwvj1UexG3vgvPm6ttxB
j7WoFy6tbRuDSxIbySiAwB4+xd0c+saIJpISP0+kAjT+ytfm6SZrA72WdEssY57Het8b4uhpRFCZJ8RH0gIL7QpJzuqvwwHUzVlz1AhLkcCPtagXLq1tG4NLEhvJKIDA
SmE0Q4DFQSR3jZb1WDWJfT8Hru8QkGKOMRYVDyLTQwTS/z352BNDdzmNYEwVR5/YYe3DnIpseeNc+xiGgCRH6a2TuLiRTboQXOaBad9FM5t39eJn8Uhh7WNDUfm7Zgrz
5y+lHQbUbWrdEx3ck1ijKo+1qBcurW0bg0sSG8kogMAhHCnLaSKqTsaFOkZn5IKDbgIsZ/OQODko6hQVsjDpd9/X329WjS8kG0eS/Uz5cImPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwOCABLjGX+83ZJjUdyx0FNvbLBOP9Pzd1AG6qUEjyql37PSJD67dlHkxZ5qJ70R+P3OD9pDjR4KrJBrEEaOfccWPtagXLq1tG4NLEhvJKIDA
8wXNLQrCkRVCQ6fSVD96z5EsV2/wLkC3/CuNN5vAQ1b9szNSM0L8NHNfAkTDNYV7bM52Edpq2Hgb3DctNgIwwKlbnXuGFUUmtV1GPME/NEACU88SnMgHnPUg1XJ+twyo
rf9pTqkh5eDvqkR6cqOb5WO1njvJVUfdph2Wm6K8vo/6ElBffe8ELvzIO1vSRDCi8af//WVDudRkGyjX+82j8Lwpvm97BH2mdJUBOY0d/150vv4ch/Gi5439gNetQ0g7
j7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAL71iCCWp2Yai5SbdqA3hwkVMM2q+NuDDLiBcXfW8riwpQMzFdJs6rRieGTCECDa2
X/wUSIn6kVuf3MS1c0URTY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAj7WoFy6tbRuDSxIbySiAwIkTtD4+JQAJdIisJ02TW4yovFIlLsru1JxXVHHindY+
rJXWXmWQM1XwNrI2nlEg72kDB+Lka186XwdmQlch/W6tfVSUwHI2FdOIbbQxC/JIj7WoFy6tbRuDSxIbySiAwI+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDA
j7WoFy6tbRuDSxIbySiAwHJak/JIchU5Hc5Ls+ruWtJm2riyWpJves/Qom6GPOb/j7WoFy6tbRuDSxIbySiAwLKDsr4oKygtbg6zqZ+nBsBcyO2qyQ5L6YzC4eV7Dvx9
OY/Hq0X/DvtVu9dBWbeCHY+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAzlokkZ3bSHowciWw+4nVP57Ef+3lvAOSv8YkLfyF7jscJlhJoHNQMCNrye9EyYNk
GixVDziA0f96l1TVhYzLyBZiqG6k/7/0iZ9W2+z4B+TlAaPdT9u726re7iWcd+fvme+sdKVX9jm7XdZs73HkdC9br6mznTtx7s4Eu+kTR8w7021YAuhU3XRSSyCitWjj
n0YxJ6y0avbPygVoMCoL7I+1qBcurW0bg0sSG8kogMCPtagXLq1tG4NLEhvJKIDAETsLCrcQ6fNtlYbORQULk9dJBVzn1WRkDKZVoVce+Fdzg/aQ40eCqyQaxBGjn3HF
j7WoFy6tbRuDSxIbySiAwLvjDjAQEB6k4KJDSerd3MrgDtsVjtRR+iGuTxghxDevm2lQRDoecMLFYzrrakyNQydCtfuGIUam17WdlqxVEZCPtagXLq1tG4NLEhvJKIDA
soOyvigrKC1uDrOpn6cGwFpAMziTBHOrnUuONdgaBT03EDGiCLj9ZFT0AIX0IQ9h9hMo5HCkK5/RMwWxkN/UFqaBEikicyj6zVQrJkuR1n/jMe/3Mb0/N7MEzxOFNODH
W74LjjSPM8i8zaVfYVyauicmyIGfdK6q5dloUYhNgHePal/ccQmjcnsBywQ9NAFHqVude4YVRSa1XUY8wT80QGK/rScqFJ3DoZa4wCDR29Yl0TF+yuCPf3JG1rzh1B5B
bfLA1EcB/Hwhbqd71DLez/etSo46JNIh2FMgyDkdWK5bPD4L3F6POR0TK26EOwPafG0MHAtlJQeTc5ESrnFVpZx+7e+P4eF0qz8myC/v7y3IKDQRTJPxz6vWZ+IlR0jQ
Gtd/3Ce2xs2Z+SKr6NJ+cRCAA1WdpGdHH8EMgS7yr4+g96O5ZNtO+Zr0ePRhXDnpHYIzagPvprLvLXRmsKjPeLw08eYqNONu7zSbqlNYw5Nc87IOTcgLSaToZt+lYHjU
s4m5tMwJf9i3Bw06+dMY1qOVdyR65Qg15/FcUH7chZpGTprZInZ7ICLjXI+/0RJtT9/3tgUcUYLbigmL1XSrHzG6mHHxa6dS++mMcrWoh1SX9hHM3b2TRIX+ePSz5afN
KRINuworNlbrQ1twv+fa7zDzj/DzbcN9JHYk//LF6ozn0T6JX3dWElj1KtFzrmU+/wCw8Z9KwwNpYlpQeXe/v8LEG8gzkH7pa8+RHDbOuac5IocDABHZ274kbp3zjv1g
iWAtes8YLIyPCQyyEKubni72MfLL266b6+sgpJanfnnCeUdRCGwlm/hK7BEEPoMKbfLA1EcB/Hwhbqd71DLez/etSo46JNIh2FMgyDkdWK7TpOxHkPPEz965i0+DpF64
xikIRr4+YY6/wCwuDy/AkEN5baQkSHB9pOEoOmjqlyX8CvFL9nXrqXZvAioIb0/7a3luoiFeVzf2kj6Xu+ek64637zgO76y0hrqTgEkMsp7ocD3FVfM9fk3LC40CFkF3
M+a96Sq5yv4QLhj9edYASWGL0ViS/C2p2MQ/nlIRTFJDzXA+Co2wAXim1Hl8HV3qqLxSJS7K7tScV1Rx4p3WPqyV1l5lkDNV8DayNp5RIO/C3W6hHB5TQgyrroVR1uZU
c9HLp9/sCSBW/fpDsayVouGfAZkK8y5pWcW1fY069HpzLrjLT8eGegXH3zYexSfQPFOxW5sBxqpzoQ62LQrkCHfDmf8g8eT6reZZ0SMjSpHOY9UtXASwPn/UAjz+FmAW
fqUB0kR2LGEPLXWgcs7Uqa95HHg9XwAbrkcdIWcLng2ccOiE6vsYYXZIEKChAChWC/t9UQmtKSinlPAi4FMyohgZeUPmY+NzxQ1kv6WUZFpdOBL2/fUR/5ffK37RzKIw
aguS2poQU5M4DZKzQigO8F3/QGU2g9KB+ebd4MtyCLNQwT1qwumgy/xwcp16fn6TEN5qeuVaiuvil4v7TmNH4nl6yzhVLlcXtxiohkB0h/NoOBVgFym0YmMyEI2taIsM
MdpFCL12+/28jP+enpyzz7Pqzge+g22Bp+dJaQJvBsAG7KhKXaNRzDDKbHEZdUIxv6kGvStasWk6bchf4439nX9V8AW63PFScoHTEBs/EB3hk5FfpJ30+nR+e2AXhc43
rER3u6YLpBHdoDJFV8jk/kgiNMmlLyBvITmWm1xTxPub0p1ntPYPZfN1S4p9pZq7MXelSorXtr3zdFgo3nwtaIjglaOBhD39Q55l67yPFarDGGA1khQJj80wFpiA8Klj
nRu+6k9KS/9uQT10PQ6gctmrUwMSdToDkD4QIDzcjdz/J3HNm5S9KM0akq9RtYkKWKIz9Q9vwx4R442Tc3bJr/v67fpar9+Ur4kyC8f12riuHGZmTOMKp5WBTPlxD5Rn
EzwknVvQhcfrCyDyf7FsNZx+7e+P4eF0qz8myC/v7y0Tii995Gdy1GBO045+WeTvLeI6pGZtq4zwHnQkAHmYtPtuOwoRIlDbrU6kkB+YdXg0K+yo1olyeZNhtpcCFHyP
ZeSrJrsoSzXeAafPFoq72+P0540tlxjkEundPIzBqIhSfVH91YqlBpKeRcKkUwngi+/7Sx1D0hFJIh7QwFSXe7Pqzge+g22Bp+dJaQJvBsDZ48vSGPe50jeZqqnsx5Ab
Vmy/r8r/TW80TSVz1xmdNE+w5QjoOrBFzwjKa0tqg8LGAqv/JMqZONnPGH74C1FB/jvL+whHBap4wXXMmC/dxSZXBueQzzuu3gEjEpRhvfuIT2lXUm7tMDSanzkHJkfL
nYAecz8wEyy01fVEpd7p7sMYYDWSFAmPzTAWmIDwqWN+AHLHs3XE9AiRBQLd5q3OE4smA+4BlMXGETyZEPyIn0zKYYQsWND4dn/FfHVSVSZSzqqTvA5kf+1gOMwbM8lH
+HzK+ij0uRU489FhKHr+7X9V8AW63PFScoHTEBs/EB2oGBQaPNZ6v/RB6+PGwoT6sxjSsOKDN55jl2DXhsBmD4qeDlJ+YMPjdTyCMtZq1jPhPHbc0qCa9cidluxSNRPR
WzXU3PazDsKyEoFITyPF6gGTgzoMjaMtfQckVs+jeJVuCR73WopvhmiAf+KHLwqZgsy6dg4kKSCoDf8fYe5pzFEvNWUmHx7uJI8uQROazSkJRy3Ki5LKaHQh1ruFfPGl
0oOK1x8LJ436PozPxcMJgZy/pF/0HjYgIFz0hTluMNS/meV+kuy3KCyDfk7PVohmN6PO0HcqD+6PaWOKB/XyE3mgPTnDdFOqrPjVWXFRRECgVQsi5yjZvUhhT5ynLTpM
wLSiyrUR8/8AlitblUypSpx+7e+P4eF0qz8myC/v7y3I5ynYRc1qSW5AhibDiFcW93TGv9Z4p+sxso7At3kNW2Ju4OJ43r/pgsYnaHd3zJK4MzW5VXwenbkHwD3pkHgc
/Pn880DGdrDRslsmbaOY4ogo5nqny+DmDItt9IwXS9lY74SCvxNPJYvCrt3kDo9dqxjKnYE3mA4ut7WtibPzcByOGwwQaWWx1VHN8+kKrptYojP1D2/DHhHjjZNzdsmv
UR0vPAY7/cEcGPsyeZPoyehwPcVV8z1+TcsLjQIWQXcTT4BfvGL9/v/V3Rj9VtkOwEBwuPTrmsXmyWZFoZu3a8HGjQWiLqDKhGWbZRRAsTMafSyOxdjsup0BGSi2/OU/
L7d1xjVa3ojtrXnCmMwkuJ0bvupPSkv/bkE9dD0OoHL3rUqOOiTSIdhTIMg5HViuzQOQSv3Ql7f3vzjpm8oYf/MwmexKfF4fsPv8rjrSS+3dxvKh9ZMhw/36feIv7oOk
abyi7UxFF8IqLh9pPqc3yRz9PCTH5YJ7vPRanAPomj8xi1iGOXcwrc5LhPeQnCfdrhTm8EqyrFAh0eisT/jjK7p179MSB44+j9nNm5E9m5CEhHek0+xn+ThfPlffoOs1
dcvfuaqMep524XAvNLI1Puy9jfkulbOK3m4jT1/Vel1Hwg5VCMOD6FFLp/nDSoqdCRLqDKaHHciNZeLDCImGu/uVToQDN7l6VTgJ7d1zHDrwhkp+UMkvKGZ0UVnOJcJQ
d8uXi0x7jTiy03xlTmIsGJ/HP+B5nem8KqMimrOZM+UIFDXUoORH6Kd7xifjxxPVLY0qbdm0OXhuREFeDj/CPdZOfMcylxrg6WxIqxkwbg5wnFrhurYcHg6JOPpNCKsG
HHnT41v1f1YjpgTjLbF13THaRQi9dvv9vIz/np6cs8+z6s4HvoNtgafnSWkCbwbABuyoSl2jUcwwymxxGXVCMcMyVVNlVj64AEyLm2HQFeapW517hhVFJrVdRjzBPzRA
0308cxY9VZeH1+nozoAA7GHyX3w9WDTEk+GlvhSk/cKsu1TIihdgjStH17G7//vk3t3vorCuJ45+2cFpYnv8z0qUWmlyqcA9dxlkV6/4yapd7ScA8YNNWfGqjlbe9koG
5Kwy3aY6ak4hAn+3/PWgOsMYYDWSFAmPzTAWmIDwqWOL7/tLHUPSEUkiHtDAVJd7kLLqDQTBRtnd0vjH3Mk1TqlbnXuGFUUmtV1GPME/NEAqHwEogofTV+r+Pg6rjObk
An8mSUsVqiYI37xmV58LtK8zmuSt2Q0hf0ISONNcl700K+yo1olyeZNhtpcCFHyPCObB8riFBrJSzQ/3Y/Qxqn2kCjSsFgKj6D7HNrGHAPiaIj3frYsws81ln2baUsNG
BWsYpleyjclbwUrkJJzjnhLJscF3QF5S9Tc1gT6HWFxMQjguUouKUXwfQ/28qrFUJZZ7tiHGdBzrp5cU6RkUn9logjS8qNH7U6Rwect+NiL/ALDxn0rDA2liWlB5d7+/
i+/7Sx1D0hFJIh7QwFSXe7Pqzge+g22Bp+dJaQJvBsDZ48vSGPe50jeZqqnsx5AbxMAWKjsY4s1ykAcWBq2l2CMCmFgSqI5hOZKzPA8htzmj/wR8LAsOPLIpR7ge0I/U
`pragma protect end_protected
